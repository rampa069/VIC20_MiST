
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"44",x"6c",x"38",x"10"),
     1 => (x"bc",x"1c",x"00",x"00"),
     2 => (x"1c",x"3c",x"60",x"e0"),
     3 => (x"64",x"44",x"00",x"00"),
     4 => (x"44",x"4c",x"5c",x"74"),
     5 => (x"08",x"08",x"00",x"00"),
     6 => (x"41",x"41",x"77",x"3e"),
     7 => (x"00",x"00",x"00",x"00"),
     8 => (x"00",x"00",x"7f",x"7f"),
     9 => (x"41",x"41",x"00",x"00"),
    10 => (x"08",x"08",x"3e",x"77"),
    11 => (x"01",x"01",x"02",x"00"),
    12 => (x"01",x"02",x"02",x"03"),
    13 => (x"7f",x"7f",x"7f",x"00"),
    14 => (x"7f",x"7f",x"7f",x"7f"),
    15 => (x"1c",x"08",x"08",x"00"),
    16 => (x"7f",x"3e",x"3e",x"1c"),
    17 => (x"3e",x"7f",x"7f",x"7f"),
    18 => (x"08",x"1c",x"1c",x"3e"),
    19 => (x"18",x"10",x"00",x"08"),
    20 => (x"10",x"18",x"7c",x"7c"),
    21 => (x"30",x"10",x"00",x"00"),
    22 => (x"10",x"30",x"7c",x"7c"),
    23 => (x"60",x"30",x"10",x"00"),
    24 => (x"06",x"1e",x"78",x"60"),
    25 => (x"3c",x"66",x"42",x"00"),
    26 => (x"42",x"66",x"3c",x"18"),
    27 => (x"6a",x"38",x"78",x"00"),
    28 => (x"38",x"6c",x"c6",x"c2"),
    29 => (x"00",x"00",x"60",x"00"),
    30 => (x"60",x"00",x"00",x"60"),
    31 => (x"5b",x"5e",x"0e",x"00"),
    32 => (x"1e",x"0e",x"5d",x"5c"),
    33 => (x"eb",x"c2",x"4c",x"71"),
    34 => (x"c0",x"4d",x"bf",x"d6"),
    35 => (x"74",x"1e",x"c0",x"4b"),
    36 => (x"87",x"c7",x"02",x"ab"),
    37 => (x"c0",x"48",x"a6",x"c4"),
    38 => (x"c4",x"87",x"c5",x"78"),
    39 => (x"78",x"c1",x"48",x"a6"),
    40 => (x"73",x"1e",x"66",x"c4"),
    41 => (x"87",x"df",x"ee",x"49"),
    42 => (x"e0",x"c0",x"86",x"c8"),
    43 => (x"87",x"ef",x"ef",x"49"),
    44 => (x"6a",x"4a",x"a5",x"c4"),
    45 => (x"87",x"f0",x"f0",x"49"),
    46 => (x"cb",x"87",x"c6",x"f1"),
    47 => (x"c8",x"83",x"c1",x"85"),
    48 => (x"ff",x"04",x"ab",x"b7"),
    49 => (x"26",x"26",x"87",x"c7"),
    50 => (x"26",x"4c",x"26",x"4d"),
    51 => (x"1e",x"4f",x"26",x"4b"),
    52 => (x"eb",x"c2",x"4a",x"71"),
    53 => (x"eb",x"c2",x"5a",x"da"),
    54 => (x"78",x"c7",x"48",x"da"),
    55 => (x"87",x"dd",x"fe",x"49"),
    56 => (x"73",x"1e",x"4f",x"26"),
    57 => (x"c0",x"4a",x"71",x"1e"),
    58 => (x"d3",x"03",x"aa",x"b7"),
    59 => (x"f2",x"d0",x"c2",x"87"),
    60 => (x"87",x"c4",x"05",x"bf"),
    61 => (x"87",x"c2",x"4b",x"c1"),
    62 => (x"d0",x"c2",x"4b",x"c0"),
    63 => (x"87",x"c4",x"5b",x"f6"),
    64 => (x"5a",x"f6",x"d0",x"c2"),
    65 => (x"bf",x"f2",x"d0",x"c2"),
    66 => (x"c1",x"9a",x"c1",x"4a"),
    67 => (x"ec",x"49",x"a2",x"c0"),
    68 => (x"48",x"fc",x"87",x"e8"),
    69 => (x"bf",x"f2",x"d0",x"c2"),
    70 => (x"87",x"ef",x"fe",x"78"),
    71 => (x"c4",x"4a",x"71",x"1e"),
    72 => (x"49",x"72",x"1e",x"66"),
    73 => (x"26",x"87",x"f5",x"e9"),
    74 => (x"c2",x"1e",x"4f",x"26"),
    75 => (x"49",x"bf",x"f2",x"d0"),
    76 => (x"c2",x"87",x"f3",x"e6"),
    77 => (x"e8",x"48",x"ce",x"eb"),
    78 => (x"eb",x"c2",x"78",x"bf"),
    79 => (x"bf",x"ec",x"48",x"ca"),
    80 => (x"ce",x"eb",x"c2",x"78"),
    81 => (x"c3",x"49",x"4a",x"bf"),
    82 => (x"b7",x"c8",x"99",x"ff"),
    83 => (x"71",x"48",x"72",x"2a"),
    84 => (x"d6",x"eb",x"c2",x"b0"),
    85 => (x"0e",x"4f",x"26",x"58"),
    86 => (x"5d",x"5c",x"5b",x"5e"),
    87 => (x"ff",x"4b",x"71",x"0e"),
    88 => (x"eb",x"c2",x"87",x"c8"),
    89 => (x"50",x"c0",x"48",x"c9"),
    90 => (x"d9",x"e6",x"49",x"73"),
    91 => (x"4c",x"49",x"70",x"87"),
    92 => (x"ee",x"cb",x"9c",x"c2"),
    93 => (x"87",x"c2",x"cb",x"49"),
    94 => (x"c2",x"4d",x"49",x"70"),
    95 => (x"bf",x"97",x"c9",x"eb"),
    96 => (x"87",x"e2",x"c1",x"05"),
    97 => (x"c2",x"49",x"66",x"d0"),
    98 => (x"99",x"bf",x"d2",x"eb"),
    99 => (x"d4",x"87",x"d6",x"05"),
   100 => (x"eb",x"c2",x"49",x"66"),
   101 => (x"05",x"99",x"bf",x"ca"),
   102 => (x"49",x"73",x"87",x"cb"),
   103 => (x"70",x"87",x"e7",x"e5"),
   104 => (x"c1",x"c1",x"02",x"98"),
   105 => (x"fe",x"4c",x"c1",x"87"),
   106 => (x"49",x"75",x"87",x"c0"),
   107 => (x"70",x"87",x"d7",x"ca"),
   108 => (x"87",x"c6",x"02",x"98"),
   109 => (x"48",x"c9",x"eb",x"c2"),
   110 => (x"eb",x"c2",x"50",x"c1"),
   111 => (x"05",x"bf",x"97",x"c9"),
   112 => (x"c2",x"87",x"e3",x"c0"),
   113 => (x"49",x"bf",x"d2",x"eb"),
   114 => (x"05",x"99",x"66",x"d0"),
   115 => (x"c2",x"87",x"d6",x"ff"),
   116 => (x"49",x"bf",x"ca",x"eb"),
   117 => (x"05",x"99",x"66",x"d4"),
   118 => (x"73",x"87",x"ca",x"ff"),
   119 => (x"87",x"e6",x"e4",x"49"),
   120 => (x"fe",x"05",x"98",x"70"),
   121 => (x"48",x"74",x"87",x"ff"),
   122 => (x"0e",x"87",x"dc",x"fb"),
   123 => (x"5d",x"5c",x"5b",x"5e"),
   124 => (x"c0",x"86",x"f4",x"0e"),
   125 => (x"bf",x"ec",x"4c",x"4d"),
   126 => (x"48",x"a6",x"c4",x"7e"),
   127 => (x"bf",x"d6",x"eb",x"c2"),
   128 => (x"c0",x"1e",x"c1",x"78"),
   129 => (x"fd",x"49",x"c7",x"1e"),
   130 => (x"86",x"c8",x"87",x"cd"),
   131 => (x"cd",x"02",x"98",x"70"),
   132 => (x"fb",x"49",x"ff",x"87"),
   133 => (x"da",x"c1",x"87",x"cc"),
   134 => (x"87",x"ea",x"e3",x"49"),
   135 => (x"eb",x"c2",x"4d",x"c1"),
   136 => (x"02",x"bf",x"97",x"c9"),
   137 => (x"d2",x"cd",x"87",x"c3"),
   138 => (x"ce",x"eb",x"c2",x"87"),
   139 => (x"d0",x"c2",x"4b",x"bf"),
   140 => (x"c0",x"05",x"bf",x"f2"),
   141 => (x"fd",x"c3",x"87",x"e9"),
   142 => (x"87",x"ca",x"e3",x"49"),
   143 => (x"e3",x"49",x"fa",x"c3"),
   144 => (x"49",x"73",x"87",x"c4"),
   145 => (x"71",x"99",x"ff",x"c3"),
   146 => (x"fb",x"49",x"c0",x"1e"),
   147 => (x"49",x"73",x"87",x"ce"),
   148 => (x"71",x"29",x"b7",x"c8"),
   149 => (x"fb",x"49",x"c1",x"1e"),
   150 => (x"86",x"c8",x"87",x"c2"),
   151 => (x"c2",x"87",x"f9",x"c5"),
   152 => (x"4b",x"bf",x"d2",x"eb"),
   153 => (x"87",x"dd",x"02",x"9b"),
   154 => (x"bf",x"ee",x"d0",x"c2"),
   155 => (x"87",x"d6",x"c7",x"49"),
   156 => (x"c4",x"05",x"98",x"70"),
   157 => (x"d2",x"4b",x"c0",x"87"),
   158 => (x"49",x"e0",x"c2",x"87"),
   159 => (x"c2",x"87",x"fb",x"c6"),
   160 => (x"c6",x"58",x"f2",x"d0"),
   161 => (x"ee",x"d0",x"c2",x"87"),
   162 => (x"73",x"78",x"c0",x"48"),
   163 => (x"05",x"99",x"c2",x"49"),
   164 => (x"eb",x"c3",x"87",x"cd"),
   165 => (x"87",x"ee",x"e1",x"49"),
   166 => (x"99",x"c2",x"49",x"70"),
   167 => (x"fb",x"87",x"c2",x"02"),
   168 => (x"c1",x"49",x"73",x"4c"),
   169 => (x"87",x"cd",x"05",x"99"),
   170 => (x"e1",x"49",x"f4",x"c3"),
   171 => (x"49",x"70",x"87",x"d8"),
   172 => (x"c2",x"02",x"99",x"c2"),
   173 => (x"73",x"4c",x"fa",x"87"),
   174 => (x"05",x"99",x"c8",x"49"),
   175 => (x"f5",x"c3",x"87",x"cd"),
   176 => (x"87",x"c2",x"e1",x"49"),
   177 => (x"99",x"c2",x"49",x"70"),
   178 => (x"c2",x"87",x"d4",x"02"),
   179 => (x"02",x"bf",x"da",x"eb"),
   180 => (x"c1",x"48",x"87",x"c9"),
   181 => (x"de",x"eb",x"c2",x"88"),
   182 => (x"ff",x"87",x"c2",x"58"),
   183 => (x"73",x"4d",x"c1",x"4c"),
   184 => (x"05",x"99",x"c4",x"49"),
   185 => (x"f2",x"c3",x"87",x"cd"),
   186 => (x"87",x"da",x"e0",x"49"),
   187 => (x"99",x"c2",x"49",x"70"),
   188 => (x"c2",x"87",x"db",x"02"),
   189 => (x"7e",x"bf",x"da",x"eb"),
   190 => (x"a8",x"b7",x"c7",x"48"),
   191 => (x"6e",x"87",x"cb",x"03"),
   192 => (x"c2",x"80",x"c1",x"48"),
   193 => (x"c0",x"58",x"de",x"eb"),
   194 => (x"4c",x"fe",x"87",x"c2"),
   195 => (x"fd",x"c3",x"4d",x"c1"),
   196 => (x"f1",x"df",x"ff",x"49"),
   197 => (x"c2",x"49",x"70",x"87"),
   198 => (x"87",x"d5",x"02",x"99"),
   199 => (x"bf",x"da",x"eb",x"c2"),
   200 => (x"87",x"c9",x"c0",x"02"),
   201 => (x"48",x"da",x"eb",x"c2"),
   202 => (x"c2",x"c0",x"78",x"c0"),
   203 => (x"c1",x"4c",x"fd",x"87"),
   204 => (x"49",x"fa",x"c3",x"4d"),
   205 => (x"87",x"ce",x"df",x"ff"),
   206 => (x"99",x"c2",x"49",x"70"),
   207 => (x"c2",x"87",x"d9",x"02"),
   208 => (x"48",x"bf",x"da",x"eb"),
   209 => (x"03",x"a8",x"b7",x"c7"),
   210 => (x"c2",x"87",x"c9",x"c0"),
   211 => (x"c7",x"48",x"da",x"eb"),
   212 => (x"87",x"c2",x"c0",x"78"),
   213 => (x"4d",x"c1",x"4c",x"fc"),
   214 => (x"03",x"ac",x"b7",x"c0"),
   215 => (x"c4",x"87",x"d1",x"c0"),
   216 => (x"d8",x"c1",x"4a",x"66"),
   217 => (x"c0",x"02",x"6a",x"82"),
   218 => (x"4b",x"6a",x"87",x"c6"),
   219 => (x"0f",x"73",x"49",x"74"),
   220 => (x"f0",x"c3",x"1e",x"c0"),
   221 => (x"49",x"da",x"c1",x"1e"),
   222 => (x"c8",x"87",x"dc",x"f7"),
   223 => (x"02",x"98",x"70",x"86"),
   224 => (x"c8",x"87",x"e2",x"c0"),
   225 => (x"eb",x"c2",x"48",x"a6"),
   226 => (x"c8",x"78",x"bf",x"da"),
   227 => (x"91",x"cb",x"49",x"66"),
   228 => (x"71",x"48",x"66",x"c4"),
   229 => (x"6e",x"7e",x"70",x"80"),
   230 => (x"c8",x"c0",x"02",x"bf"),
   231 => (x"4b",x"bf",x"6e",x"87"),
   232 => (x"73",x"49",x"66",x"c8"),
   233 => (x"02",x"9d",x"75",x"0f"),
   234 => (x"c2",x"87",x"c8",x"c0"),
   235 => (x"49",x"bf",x"da",x"eb"),
   236 => (x"c2",x"87",x"ca",x"f3"),
   237 => (x"02",x"bf",x"f6",x"d0"),
   238 => (x"49",x"87",x"dd",x"c0"),
   239 => (x"70",x"87",x"c7",x"c2"),
   240 => (x"d3",x"c0",x"02",x"98"),
   241 => (x"da",x"eb",x"c2",x"87"),
   242 => (x"f0",x"f2",x"49",x"bf"),
   243 => (x"f4",x"49",x"c0",x"87"),
   244 => (x"d0",x"c2",x"87",x"d0"),
   245 => (x"78",x"c0",x"48",x"f6"),
   246 => (x"ea",x"f3",x"8e",x"f4"),
   247 => (x"5b",x"5e",x"0e",x"87"),
   248 => (x"1e",x"0e",x"5d",x"5c"),
   249 => (x"eb",x"c2",x"4c",x"71"),
   250 => (x"c1",x"49",x"bf",x"d6"),
   251 => (x"c1",x"4d",x"a1",x"cd"),
   252 => (x"7e",x"69",x"81",x"d1"),
   253 => (x"cf",x"02",x"9c",x"74"),
   254 => (x"4b",x"a5",x"c4",x"87"),
   255 => (x"eb",x"c2",x"7b",x"74"),
   256 => (x"f3",x"49",x"bf",x"d6"),
   257 => (x"7b",x"6e",x"87",x"c9"),
   258 => (x"c4",x"05",x"9c",x"74"),
   259 => (x"c2",x"4b",x"c0",x"87"),
   260 => (x"73",x"4b",x"c1",x"87"),
   261 => (x"87",x"ca",x"f3",x"49"),
   262 => (x"c7",x"02",x"66",x"d4"),
   263 => (x"87",x"da",x"49",x"87"),
   264 => (x"87",x"c2",x"4a",x"70"),
   265 => (x"d0",x"c2",x"4a",x"c0"),
   266 => (x"f2",x"26",x"5a",x"fa"),
   267 => (x"00",x"00",x"87",x"d9"),
   268 => (x"00",x"00",x"00",x"00"),
   269 => (x"00",x"00",x"00",x"00"),
   270 => (x"71",x"1e",x"00",x"00"),
   271 => (x"bf",x"c8",x"ff",x"4a"),
   272 => (x"48",x"a1",x"72",x"49"),
   273 => (x"ff",x"1e",x"4f",x"26"),
   274 => (x"fe",x"89",x"bf",x"c8"),
   275 => (x"c0",x"c0",x"c0",x"c0"),
   276 => (x"c4",x"01",x"a9",x"c0"),
   277 => (x"c2",x"4a",x"c0",x"87"),
   278 => (x"72",x"4a",x"c1",x"87"),
   279 => (x"0e",x"4f",x"26",x"48"),
   280 => (x"5d",x"5c",x"5b",x"5e"),
   281 => (x"7e",x"71",x"1e",x"0e"),
   282 => (x"6e",x"4b",x"d4",x"ff"),
   283 => (x"de",x"eb",x"c2",x"1e"),
   284 => (x"d8",x"cf",x"fe",x"49"),
   285 => (x"70",x"86",x"c4",x"87"),
   286 => (x"c3",x"02",x"9d",x"4d"),
   287 => (x"eb",x"c2",x"87",x"c3"),
   288 => (x"6e",x"4c",x"bf",x"e6"),
   289 => (x"d0",x"e2",x"fe",x"49"),
   290 => (x"48",x"d0",x"ff",x"87"),
   291 => (x"c1",x"78",x"c5",x"c8"),
   292 => (x"4a",x"c0",x"7b",x"d6"),
   293 => (x"82",x"c1",x"7b",x"15"),
   294 => (x"aa",x"b7",x"e0",x"c0"),
   295 => (x"ff",x"87",x"f5",x"04"),
   296 => (x"78",x"c4",x"48",x"d0"),
   297 => (x"c1",x"78",x"c5",x"c8"),
   298 => (x"7b",x"c1",x"7b",x"d3"),
   299 => (x"9c",x"74",x"78",x"c4"),
   300 => (x"87",x"fc",x"c1",x"02"),
   301 => (x"7e",x"ce",x"da",x"c2"),
   302 => (x"8c",x"4d",x"c0",x"c8"),
   303 => (x"03",x"ac",x"b7",x"c0"),
   304 => (x"c0",x"c8",x"87",x"c6"),
   305 => (x"4c",x"c0",x"4d",x"a4"),
   306 => (x"97",x"ff",x"e6",x"c2"),
   307 => (x"99",x"d0",x"49",x"bf"),
   308 => (x"c0",x"87",x"d2",x"02"),
   309 => (x"de",x"eb",x"c2",x"1e"),
   310 => (x"cc",x"d1",x"fe",x"49"),
   311 => (x"70",x"86",x"c4",x"87"),
   312 => (x"ef",x"c0",x"4a",x"49"),
   313 => (x"ce",x"da",x"c2",x"87"),
   314 => (x"de",x"eb",x"c2",x"1e"),
   315 => (x"f8",x"d0",x"fe",x"49"),
   316 => (x"70",x"86",x"c4",x"87"),
   317 => (x"d0",x"ff",x"4a",x"49"),
   318 => (x"78",x"c5",x"c8",x"48"),
   319 => (x"6e",x"7b",x"d4",x"c1"),
   320 => (x"6e",x"7b",x"bf",x"97"),
   321 => (x"70",x"80",x"c1",x"48"),
   322 => (x"05",x"8d",x"c1",x"7e"),
   323 => (x"ff",x"87",x"f0",x"ff"),
   324 => (x"78",x"c4",x"48",x"d0"),
   325 => (x"c5",x"05",x"9a",x"72"),
   326 => (x"c0",x"48",x"c0",x"87"),
   327 => (x"1e",x"c1",x"87",x"e5"),
   328 => (x"49",x"de",x"eb",x"c2"),
   329 => (x"87",x"e0",x"ce",x"fe"),
   330 => (x"9c",x"74",x"86",x"c4"),
   331 => (x"87",x"c4",x"fe",x"05"),
   332 => (x"c8",x"48",x"d0",x"ff"),
   333 => (x"d3",x"c1",x"78",x"c5"),
   334 => (x"c4",x"7b",x"c0",x"7b"),
   335 => (x"c2",x"48",x"c1",x"78"),
   336 => (x"26",x"48",x"c0",x"87"),
   337 => (x"4c",x"26",x"4d",x"26"),
   338 => (x"4f",x"26",x"4b",x"26"),
   339 => (x"71",x"1e",x"73",x"1e"),
   340 => (x"02",x"66",x"c8",x"4a"),
   341 => (x"c1",x"4b",x"87",x"ce"),
   342 => (x"ce",x"02",x"8b",x"d3"),
   343 => (x"02",x"8b",x"c1",x"87"),
   344 => (x"87",x"d3",x"87",x"d0"),
   345 => (x"f6",x"fb",x"49",x"72"),
   346 => (x"72",x"87",x"cc",x"87"),
   347 => (x"87",x"ca",x"c2",x"49"),
   348 => (x"49",x"72",x"87",x"c5"),
   349 => (x"ff",x"87",x"f6",x"c2"),
   350 => (x"1e",x"00",x"87",x"ce"),
   351 => (x"bf",x"e2",x"d9",x"c2"),
   352 => (x"c2",x"b9",x"c1",x"49"),
   353 => (x"ff",x"59",x"e6",x"d9"),
   354 => (x"ff",x"c3",x"48",x"d4"),
   355 => (x"48",x"d0",x"ff",x"78"),
   356 => (x"ff",x"78",x"e1",x"c8"),
   357 => (x"78",x"c1",x"48",x"d4"),
   358 => (x"78",x"71",x"31",x"c4"),
   359 => (x"c0",x"48",x"d0",x"ff"),
   360 => (x"4f",x"26",x"78",x"e0"),
   361 => (x"fd",x"d6",x"c2",x"1e"),
   362 => (x"de",x"eb",x"c2",x"1e"),
   363 => (x"dc",x"ca",x"fe",x"49"),
   364 => (x"70",x"86",x"c4",x"87"),
   365 => (x"87",x"c3",x"02",x"98"),
   366 => (x"26",x"87",x"c0",x"ff"),
   367 => (x"4b",x"35",x"31",x"4f"),
   368 => (x"20",x"20",x"5a",x"48"),
   369 => (x"47",x"46",x"43",x"20"),
   370 => (x"4a",x"71",x"1e",x"00"),
   371 => (x"c2",x"49",x"a2",x"c4"),
   372 => (x"6a",x"48",x"f5",x"ea"),
   373 => (x"c1",x"49",x"69",x"78"),
   374 => (x"e6",x"d9",x"c2",x"b9"),
   375 => (x"87",x"db",x"fe",x"59"),
   376 => (x"87",x"d9",x"d7",x"ff"),
   377 => (x"4f",x"26",x"48",x"c1"),
   378 => (x"c4",x"4a",x"71",x"1e"),
   379 => (x"ea",x"c2",x"49",x"a2"),
   380 => (x"c2",x"7a",x"bf",x"f5"),
   381 => (x"79",x"bf",x"e2",x"d9"),
   382 => (x"71",x"1e",x"4f",x"26"),
   383 => (x"eb",x"c2",x"1e",x"4a"),
   384 => (x"c9",x"fe",x"49",x"de"),
   385 => (x"86",x"c4",x"87",x"c7"),
   386 => (x"dc",x"02",x"98",x"70"),
   387 => (x"ce",x"da",x"c2",x"87"),
   388 => (x"de",x"eb",x"c2",x"1e"),
   389 => (x"d0",x"cc",x"fe",x"49"),
   390 => (x"70",x"86",x"c4",x"87"),
   391 => (x"87",x"c9",x"02",x"98"),
   392 => (x"49",x"ce",x"da",x"c2"),
   393 => (x"c2",x"87",x"e2",x"fe"),
   394 => (x"26",x"48",x"c0",x"87"),
   395 => (x"4a",x"71",x"1e",x"4f"),
   396 => (x"de",x"eb",x"c2",x"1e"),
   397 => (x"d4",x"c8",x"fe",x"49"),
   398 => (x"70",x"86",x"c4",x"87"),
   399 => (x"87",x"de",x"02",x"98"),
   400 => (x"49",x"ce",x"da",x"c2"),
   401 => (x"c2",x"87",x"e1",x"fe"),
   402 => (x"c2",x"1e",x"ce",x"da"),
   403 => (x"fe",x"49",x"de",x"eb"),
   404 => (x"c4",x"87",x"d9",x"cc"),
   405 => (x"02",x"98",x"70",x"86"),
   406 => (x"48",x"c1",x"87",x"c4"),
   407 => (x"48",x"c0",x"87",x"c2"),
   408 => (x"00",x"00",x"4f",x"26"),
   409 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

