
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f4",x"eb",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"f4",x"eb",x"c2"),
    14 => (x"48",x"e8",x"d9",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e0",x"de"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"11",x"1e",x"4f"),
    50 => (x"78",x"08",x"d4",x"ff"),
    51 => (x"c1",x"48",x"66",x"c4"),
    52 => (x"58",x"a6",x"c8",x"88"),
    53 => (x"ed",x"05",x"98",x"70"),
    54 => (x"1e",x"4f",x"26",x"87"),
    55 => (x"c3",x"48",x"d4",x"ff"),
    56 => (x"51",x"68",x"78",x"ff"),
    57 => (x"c1",x"48",x"66",x"c4"),
    58 => (x"58",x"a6",x"c8",x"88"),
    59 => (x"eb",x"05",x"98",x"70"),
    60 => (x"1e",x"4f",x"26",x"87"),
    61 => (x"d4",x"ff",x"1e",x"73"),
    62 => (x"7b",x"ff",x"c3",x"4b"),
    63 => (x"ff",x"c3",x"4a",x"6b"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"c3",x"b1",x"72",x"32"),
    66 => (x"4a",x"6b",x"7b",x"ff"),
    67 => (x"b2",x"71",x"31",x"c8"),
    68 => (x"6b",x"7b",x"ff",x"c3"),
    69 => (x"72",x"32",x"c8",x"49"),
    70 => (x"c4",x"48",x"71",x"b1"),
    71 => (x"26",x"4d",x"26",x"87"),
    72 => (x"26",x"4b",x"26",x"4c"),
    73 => (x"5b",x"5e",x"0e",x"4f"),
    74 => (x"71",x"0e",x"5d",x"5c"),
    75 => (x"4c",x"d4",x"ff",x"4a"),
    76 => (x"ff",x"c3",x"49",x"72"),
    77 => (x"c2",x"7c",x"71",x"99"),
    78 => (x"05",x"bf",x"e8",x"d9"),
    79 => (x"66",x"d0",x"87",x"c8"),
    80 => (x"d4",x"30",x"c9",x"48"),
    81 => (x"66",x"d0",x"58",x"a6"),
    82 => (x"c3",x"29",x"d8",x"49"),
    83 => (x"7c",x"71",x"99",x"ff"),
    84 => (x"d0",x"49",x"66",x"d0"),
    85 => (x"99",x"ff",x"c3",x"29"),
    86 => (x"66",x"d0",x"7c",x"71"),
    87 => (x"c3",x"29",x"c8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"c3",x"49",x"66",x"d0"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"29",x"d0",x"49",x"72"),
    92 => (x"71",x"99",x"ff",x"c3"),
    93 => (x"c9",x"4b",x"6c",x"7c"),
    94 => (x"c3",x"4d",x"ff",x"f0"),
    95 => (x"d0",x"05",x"ab",x"ff"),
    96 => (x"7c",x"ff",x"c3",x"87"),
    97 => (x"8d",x"c1",x"4b",x"6c"),
    98 => (x"c3",x"87",x"c6",x"02"),
    99 => (x"f0",x"02",x"ab",x"ff"),
   100 => (x"fe",x"48",x"73",x"87"),
   101 => (x"c0",x"1e",x"87",x"c7"),
   102 => (x"48",x"d4",x"ff",x"49"),
   103 => (x"c1",x"78",x"ff",x"c3"),
   104 => (x"b7",x"c8",x"c3",x"81"),
   105 => (x"87",x"f1",x"04",x"a9"),
   106 => (x"73",x"1e",x"4f",x"26"),
   107 => (x"c4",x"87",x"e7",x"1e"),
   108 => (x"c0",x"4b",x"df",x"f8"),
   109 => (x"f0",x"ff",x"c0",x"1e"),
   110 => (x"fd",x"49",x"f7",x"c1"),
   111 => (x"86",x"c4",x"87",x"e7"),
   112 => (x"c0",x"05",x"a8",x"c1"),
   113 => (x"d4",x"ff",x"87",x"ea"),
   114 => (x"78",x"ff",x"c3",x"48"),
   115 => (x"c0",x"c0",x"c0",x"c1"),
   116 => (x"c0",x"1e",x"c0",x"c0"),
   117 => (x"e9",x"c1",x"f0",x"e1"),
   118 => (x"87",x"c9",x"fd",x"49"),
   119 => (x"98",x"70",x"86",x"c4"),
   120 => (x"ff",x"87",x"ca",x"05"),
   121 => (x"ff",x"c3",x"48",x"d4"),
   122 => (x"cb",x"48",x"c1",x"78"),
   123 => (x"87",x"e6",x"fe",x"87"),
   124 => (x"fe",x"05",x"8b",x"c1"),
   125 => (x"48",x"c0",x"87",x"fd"),
   126 => (x"1e",x"87",x"e6",x"fc"),
   127 => (x"d4",x"ff",x"1e",x"73"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"1e",x"c0",x"4b",x"d3"),
   130 => (x"c1",x"f0",x"ff",x"c0"),
   131 => (x"d4",x"fc",x"49",x"c1"),
   132 => (x"70",x"86",x"c4",x"87"),
   133 => (x"87",x"ca",x"05",x"98"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"48",x"c1",x"78",x"ff"),
   136 => (x"f1",x"fd",x"87",x"cb"),
   137 => (x"05",x"8b",x"c1",x"87"),
   138 => (x"c0",x"87",x"db",x"ff"),
   139 => (x"87",x"f1",x"fb",x"48"),
   140 => (x"5c",x"5b",x"5e",x"0e"),
   141 => (x"4c",x"d4",x"ff",x"0e"),
   142 => (x"c6",x"87",x"db",x"fd"),
   143 => (x"e1",x"c0",x"1e",x"ea"),
   144 => (x"49",x"c8",x"c1",x"f0"),
   145 => (x"c4",x"87",x"de",x"fb"),
   146 => (x"02",x"a8",x"c1",x"86"),
   147 => (x"ea",x"fe",x"87",x"c8"),
   148 => (x"c1",x"48",x"c0",x"87"),
   149 => (x"da",x"fa",x"87",x"e2"),
   150 => (x"cf",x"49",x"70",x"87"),
   151 => (x"c6",x"99",x"ff",x"ff"),
   152 => (x"c8",x"02",x"a9",x"ea"),
   153 => (x"87",x"d3",x"fe",x"87"),
   154 => (x"cb",x"c1",x"48",x"c0"),
   155 => (x"7c",x"ff",x"c3",x"87"),
   156 => (x"fc",x"4b",x"f1",x"c0"),
   157 => (x"98",x"70",x"87",x"f4"),
   158 => (x"87",x"eb",x"c0",x"02"),
   159 => (x"ff",x"c0",x"1e",x"c0"),
   160 => (x"49",x"fa",x"c1",x"f0"),
   161 => (x"c4",x"87",x"de",x"fa"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"ff",x"c3",x"87",x"d9"),
   164 => (x"c3",x"49",x"6c",x"7c"),
   165 => (x"7c",x"7c",x"7c",x"ff"),
   166 => (x"99",x"c0",x"c1",x"7c"),
   167 => (x"c1",x"87",x"c4",x"02"),
   168 => (x"c0",x"87",x"d5",x"48"),
   169 => (x"c2",x"87",x"d1",x"48"),
   170 => (x"87",x"c4",x"05",x"ab"),
   171 => (x"87",x"c8",x"48",x"c0"),
   172 => (x"fe",x"05",x"8b",x"c1"),
   173 => (x"48",x"c0",x"87",x"fd"),
   174 => (x"1e",x"87",x"e4",x"f9"),
   175 => (x"d9",x"c2",x"1e",x"73"),
   176 => (x"78",x"c1",x"48",x"e8"),
   177 => (x"d0",x"ff",x"4b",x"c7"),
   178 => (x"fb",x"78",x"c2",x"48"),
   179 => (x"d0",x"ff",x"87",x"c8"),
   180 => (x"c0",x"78",x"c3",x"48"),
   181 => (x"d0",x"e5",x"c0",x"1e"),
   182 => (x"f9",x"49",x"c0",x"c1"),
   183 => (x"86",x"c4",x"87",x"c7"),
   184 => (x"c1",x"05",x"a8",x"c1"),
   185 => (x"ab",x"c2",x"4b",x"87"),
   186 => (x"c0",x"87",x"c5",x"05"),
   187 => (x"87",x"f9",x"c0",x"48"),
   188 => (x"ff",x"05",x"8b",x"c1"),
   189 => (x"f7",x"fc",x"87",x"d0"),
   190 => (x"ec",x"d9",x"c2",x"87"),
   191 => (x"05",x"98",x"70",x"58"),
   192 => (x"1e",x"c1",x"87",x"cd"),
   193 => (x"c1",x"f0",x"ff",x"c0"),
   194 => (x"d8",x"f8",x"49",x"d0"),
   195 => (x"ff",x"86",x"c4",x"87"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"87",x"e0",x"c4",x"78"),
   198 => (x"58",x"f0",x"d9",x"c2"),
   199 => (x"c2",x"48",x"d0",x"ff"),
   200 => (x"48",x"d4",x"ff",x"78"),
   201 => (x"c1",x"78",x"ff",x"c3"),
   202 => (x"87",x"f5",x"f7",x"48"),
   203 => (x"5c",x"5b",x"5e",x"0e"),
   204 => (x"4a",x"71",x"0e",x"5d"),
   205 => (x"ff",x"4d",x"ff",x"c3"),
   206 => (x"7c",x"75",x"4c",x"d4"),
   207 => (x"c4",x"48",x"d0",x"ff"),
   208 => (x"7c",x"75",x"78",x"c3"),
   209 => (x"ff",x"c0",x"1e",x"72"),
   210 => (x"49",x"d8",x"c1",x"f0"),
   211 => (x"c4",x"87",x"d6",x"f7"),
   212 => (x"02",x"98",x"70",x"86"),
   213 => (x"48",x"c0",x"87",x"c5"),
   214 => (x"75",x"87",x"f0",x"c0"),
   215 => (x"7c",x"fe",x"c3",x"7c"),
   216 => (x"d4",x"1e",x"c0",x"c8"),
   217 => (x"dc",x"f5",x"49",x"66"),
   218 => (x"75",x"86",x"c4",x"87"),
   219 => (x"75",x"7c",x"75",x"7c"),
   220 => (x"e0",x"da",x"d8",x"7c"),
   221 => (x"6c",x"7c",x"75",x"4b"),
   222 => (x"c5",x"05",x"99",x"49"),
   223 => (x"05",x"8b",x"c1",x"87"),
   224 => (x"7c",x"75",x"87",x"f3"),
   225 => (x"c2",x"48",x"d0",x"ff"),
   226 => (x"f6",x"48",x"c1",x"78"),
   227 => (x"ff",x"1e",x"87",x"cf"),
   228 => (x"d0",x"ff",x"4a",x"d4"),
   229 => (x"78",x"d1",x"c4",x"48"),
   230 => (x"c1",x"7a",x"ff",x"c3"),
   231 => (x"87",x"f8",x"05",x"89"),
   232 => (x"73",x"1e",x"4f",x"26"),
   233 => (x"c5",x"4b",x"71",x"1e"),
   234 => (x"4a",x"df",x"cd",x"ee"),
   235 => (x"c3",x"48",x"d4",x"ff"),
   236 => (x"48",x"68",x"78",x"ff"),
   237 => (x"02",x"a8",x"fe",x"c3"),
   238 => (x"8a",x"c1",x"87",x"c5"),
   239 => (x"72",x"87",x"ed",x"05"),
   240 => (x"87",x"c5",x"05",x"9a"),
   241 => (x"ea",x"c0",x"48",x"c0"),
   242 => (x"02",x"9b",x"73",x"87"),
   243 => (x"66",x"c8",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c5"),
   246 => (x"66",x"c8",x"87",x"c6"),
   247 => (x"87",x"ee",x"fe",x"49"),
   248 => (x"c3",x"48",x"d4",x"ff"),
   249 => (x"73",x"78",x"78",x"ff"),
   250 => (x"87",x"c5",x"05",x"9b"),
   251 => (x"d0",x"48",x"d0",x"ff"),
   252 => (x"f4",x"48",x"c1",x"78"),
   253 => (x"73",x"1e",x"87",x"eb"),
   254 => (x"c0",x"4a",x"71",x"1e"),
   255 => (x"48",x"d4",x"ff",x"4b"),
   256 => (x"ff",x"78",x"ff",x"c3"),
   257 => (x"c3",x"c4",x"48",x"d0"),
   258 => (x"48",x"d4",x"ff",x"78"),
   259 => (x"72",x"78",x"ff",x"c3"),
   260 => (x"f0",x"ff",x"c0",x"1e"),
   261 => (x"f4",x"49",x"d1",x"c1"),
   262 => (x"86",x"c4",x"87",x"cb"),
   263 => (x"cd",x"05",x"98",x"70"),
   264 => (x"1e",x"c0",x"c8",x"87"),
   265 => (x"fd",x"49",x"66",x"cc"),
   266 => (x"86",x"c4",x"87",x"f8"),
   267 => (x"d0",x"ff",x"4b",x"70"),
   268 => (x"73",x"78",x"c2",x"48"),
   269 => (x"87",x"e9",x"f3",x"48"),
   270 => (x"5c",x"5b",x"5e",x"0e"),
   271 => (x"1e",x"c0",x"0e",x"5d"),
   272 => (x"c1",x"f0",x"ff",x"c0"),
   273 => (x"dc",x"f3",x"49",x"c9"),
   274 => (x"c2",x"1e",x"d2",x"87"),
   275 => (x"fd",x"49",x"f0",x"d9"),
   276 => (x"86",x"c8",x"87",x"d0"),
   277 => (x"84",x"c1",x"4c",x"c0"),
   278 => (x"04",x"ac",x"b7",x"d2"),
   279 => (x"d9",x"c2",x"87",x"f8"),
   280 => (x"49",x"bf",x"97",x"f0"),
   281 => (x"c1",x"99",x"c0",x"c3"),
   282 => (x"c0",x"05",x"a9",x"c0"),
   283 => (x"d9",x"c2",x"87",x"e7"),
   284 => (x"49",x"bf",x"97",x"f7"),
   285 => (x"d9",x"c2",x"31",x"d0"),
   286 => (x"4a",x"bf",x"97",x"f8"),
   287 => (x"b1",x"72",x"32",x"c8"),
   288 => (x"97",x"f9",x"d9",x"c2"),
   289 => (x"71",x"b1",x"4a",x"bf"),
   290 => (x"ff",x"ff",x"cf",x"4c"),
   291 => (x"84",x"c1",x"9c",x"ff"),
   292 => (x"e7",x"c1",x"34",x"ca"),
   293 => (x"f9",x"d9",x"c2",x"87"),
   294 => (x"c1",x"49",x"bf",x"97"),
   295 => (x"c2",x"99",x"c6",x"31"),
   296 => (x"bf",x"97",x"fa",x"d9"),
   297 => (x"2a",x"b7",x"c7",x"4a"),
   298 => (x"d9",x"c2",x"b1",x"72"),
   299 => (x"4a",x"bf",x"97",x"f5"),
   300 => (x"c2",x"9d",x"cf",x"4d"),
   301 => (x"bf",x"97",x"f6",x"d9"),
   302 => (x"ca",x"9a",x"c3",x"4a"),
   303 => (x"f7",x"d9",x"c2",x"32"),
   304 => (x"c2",x"4b",x"bf",x"97"),
   305 => (x"c2",x"b2",x"73",x"33"),
   306 => (x"bf",x"97",x"f8",x"d9"),
   307 => (x"9b",x"c0",x"c3",x"4b"),
   308 => (x"73",x"2b",x"b7",x"c6"),
   309 => (x"c1",x"81",x"c2",x"b2"),
   310 => (x"70",x"30",x"71",x"48"),
   311 => (x"75",x"48",x"c1",x"49"),
   312 => (x"72",x"4d",x"70",x"30"),
   313 => (x"71",x"84",x"c1",x"4c"),
   314 => (x"b7",x"c0",x"c8",x"94"),
   315 => (x"87",x"cc",x"06",x"ad"),
   316 => (x"2d",x"b7",x"34",x"c1"),
   317 => (x"ad",x"b7",x"c0",x"c8"),
   318 => (x"87",x"f4",x"ff",x"01"),
   319 => (x"dc",x"f0",x"48",x"74"),
   320 => (x"5b",x"5e",x"0e",x"87"),
   321 => (x"f8",x"0e",x"5d",x"5c"),
   322 => (x"d6",x"e2",x"c2",x"86"),
   323 => (x"c2",x"78",x"c0",x"48"),
   324 => (x"c0",x"1e",x"ce",x"da"),
   325 => (x"87",x"de",x"fb",x"49"),
   326 => (x"98",x"70",x"86",x"c4"),
   327 => (x"c0",x"87",x"c5",x"05"),
   328 => (x"87",x"ce",x"c9",x"48"),
   329 => (x"7e",x"c1",x"4d",x"c0"),
   330 => (x"bf",x"e4",x"f0",x"c0"),
   331 => (x"c4",x"db",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f3",x"ec"),
   334 => (x"87",x"c2",x"05",x"98"),
   335 => (x"f0",x"c0",x"7e",x"c0"),
   336 => (x"c2",x"49",x"bf",x"e0"),
   337 => (x"71",x"4a",x"e0",x"db"),
   338 => (x"dd",x"ec",x"4b",x"c8"),
   339 => (x"05",x"98",x"70",x"87"),
   340 => (x"7e",x"c0",x"87",x"c2"),
   341 => (x"fd",x"c0",x"02",x"6e"),
   342 => (x"d4",x"e1",x"c2",x"87"),
   343 => (x"e2",x"c2",x"4d",x"bf"),
   344 => (x"7e",x"bf",x"9f",x"cc"),
   345 => (x"ea",x"d6",x"c5",x"48"),
   346 => (x"87",x"c7",x"05",x"a8"),
   347 => (x"bf",x"d4",x"e1",x"c2"),
   348 => (x"6e",x"87",x"ce",x"4d"),
   349 => (x"d5",x"e9",x"ca",x"48"),
   350 => (x"87",x"c5",x"02",x"a8"),
   351 => (x"f1",x"c7",x"48",x"c0"),
   352 => (x"ce",x"da",x"c2",x"87"),
   353 => (x"f9",x"49",x"75",x"1e"),
   354 => (x"86",x"c4",x"87",x"ec"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c7",x"48",x"c0",x"87"),
   357 => (x"f0",x"c0",x"87",x"dc"),
   358 => (x"c2",x"49",x"bf",x"e0"),
   359 => (x"71",x"4a",x"e0",x"db"),
   360 => (x"c5",x"eb",x"4b",x"c8"),
   361 => (x"05",x"98",x"70",x"87"),
   362 => (x"e2",x"c2",x"87",x"c8"),
   363 => (x"78",x"c1",x"48",x"d6"),
   364 => (x"f0",x"c0",x"87",x"da"),
   365 => (x"c2",x"49",x"bf",x"e4"),
   366 => (x"71",x"4a",x"c4",x"db"),
   367 => (x"e9",x"ea",x"4b",x"c8"),
   368 => (x"02",x"98",x"70",x"87"),
   369 => (x"c0",x"87",x"c5",x"c0"),
   370 => (x"87",x"e6",x"c6",x"48"),
   371 => (x"97",x"cc",x"e2",x"c2"),
   372 => (x"d5",x"c1",x"49",x"bf"),
   373 => (x"cd",x"c0",x"05",x"a9"),
   374 => (x"cd",x"e2",x"c2",x"87"),
   375 => (x"c2",x"49",x"bf",x"97"),
   376 => (x"c0",x"02",x"a9",x"ea"),
   377 => (x"48",x"c0",x"87",x"c5"),
   378 => (x"c2",x"87",x"c7",x"c6"),
   379 => (x"bf",x"97",x"ce",x"da"),
   380 => (x"e9",x"c3",x"48",x"7e"),
   381 => (x"ce",x"c0",x"02",x"a8"),
   382 => (x"c3",x"48",x"6e",x"87"),
   383 => (x"c0",x"02",x"a8",x"eb"),
   384 => (x"48",x"c0",x"87",x"c5"),
   385 => (x"c2",x"87",x"eb",x"c5"),
   386 => (x"bf",x"97",x"d9",x"da"),
   387 => (x"c0",x"05",x"99",x"49"),
   388 => (x"da",x"c2",x"87",x"cc"),
   389 => (x"49",x"bf",x"97",x"da"),
   390 => (x"c0",x"02",x"a9",x"c2"),
   391 => (x"48",x"c0",x"87",x"c5"),
   392 => (x"c2",x"87",x"cf",x"c5"),
   393 => (x"bf",x"97",x"db",x"da"),
   394 => (x"d2",x"e2",x"c2",x"48"),
   395 => (x"48",x"4c",x"70",x"58"),
   396 => (x"e2",x"c2",x"88",x"c1"),
   397 => (x"da",x"c2",x"58",x"d6"),
   398 => (x"49",x"bf",x"97",x"dc"),
   399 => (x"da",x"c2",x"81",x"75"),
   400 => (x"4a",x"bf",x"97",x"dd"),
   401 => (x"a1",x"72",x"32",x"c8"),
   402 => (x"e3",x"e6",x"c2",x"7e"),
   403 => (x"c2",x"78",x"6e",x"48"),
   404 => (x"bf",x"97",x"de",x"da"),
   405 => (x"58",x"a6",x"c8",x"48"),
   406 => (x"bf",x"d6",x"e2",x"c2"),
   407 => (x"87",x"d4",x"c2",x"02"),
   408 => (x"bf",x"e0",x"f0",x"c0"),
   409 => (x"e0",x"db",x"c2",x"49"),
   410 => (x"4b",x"c8",x"71",x"4a"),
   411 => (x"70",x"87",x"fb",x"e7"),
   412 => (x"c5",x"c0",x"02",x"98"),
   413 => (x"c3",x"48",x"c0",x"87"),
   414 => (x"e2",x"c2",x"87",x"f8"),
   415 => (x"c2",x"4c",x"bf",x"ce"),
   416 => (x"c2",x"5c",x"f7",x"e6"),
   417 => (x"bf",x"97",x"f3",x"da"),
   418 => (x"c2",x"31",x"c8",x"49"),
   419 => (x"bf",x"97",x"f2",x"da"),
   420 => (x"c2",x"49",x"a1",x"4a"),
   421 => (x"bf",x"97",x"f4",x"da"),
   422 => (x"72",x"32",x"d0",x"4a"),
   423 => (x"da",x"c2",x"49",x"a1"),
   424 => (x"4a",x"bf",x"97",x"f5"),
   425 => (x"a1",x"72",x"32",x"d8"),
   426 => (x"91",x"66",x"c4",x"49"),
   427 => (x"bf",x"e3",x"e6",x"c2"),
   428 => (x"eb",x"e6",x"c2",x"81"),
   429 => (x"fb",x"da",x"c2",x"59"),
   430 => (x"c8",x"4a",x"bf",x"97"),
   431 => (x"fa",x"da",x"c2",x"32"),
   432 => (x"a2",x"4b",x"bf",x"97"),
   433 => (x"fc",x"da",x"c2",x"4a"),
   434 => (x"d0",x"4b",x"bf",x"97"),
   435 => (x"4a",x"a2",x"73",x"33"),
   436 => (x"97",x"fd",x"da",x"c2"),
   437 => (x"9b",x"cf",x"4b",x"bf"),
   438 => (x"a2",x"73",x"33",x"d8"),
   439 => (x"ef",x"e6",x"c2",x"4a"),
   440 => (x"eb",x"e6",x"c2",x"5a"),
   441 => (x"8a",x"c2",x"4a",x"bf"),
   442 => (x"e6",x"c2",x"92",x"74"),
   443 => (x"a1",x"72",x"48",x"ef"),
   444 => (x"87",x"ca",x"c1",x"78"),
   445 => (x"97",x"e0",x"da",x"c2"),
   446 => (x"31",x"c8",x"49",x"bf"),
   447 => (x"97",x"df",x"da",x"c2"),
   448 => (x"49",x"a1",x"4a",x"bf"),
   449 => (x"59",x"de",x"e2",x"c2"),
   450 => (x"bf",x"da",x"e2",x"c2"),
   451 => (x"c7",x"31",x"c5",x"49"),
   452 => (x"29",x"c9",x"81",x"ff"),
   453 => (x"59",x"f7",x"e6",x"c2"),
   454 => (x"97",x"e5",x"da",x"c2"),
   455 => (x"32",x"c8",x"4a",x"bf"),
   456 => (x"97",x"e4",x"da",x"c2"),
   457 => (x"4a",x"a2",x"4b",x"bf"),
   458 => (x"6e",x"92",x"66",x"c4"),
   459 => (x"f3",x"e6",x"c2",x"82"),
   460 => (x"eb",x"e6",x"c2",x"5a"),
   461 => (x"c2",x"78",x"c0",x"48"),
   462 => (x"72",x"48",x"e7",x"e6"),
   463 => (x"e6",x"c2",x"78",x"a1"),
   464 => (x"e6",x"c2",x"48",x"f7"),
   465 => (x"c2",x"78",x"bf",x"eb"),
   466 => (x"c2",x"48",x"fb",x"e6"),
   467 => (x"78",x"bf",x"ef",x"e6"),
   468 => (x"bf",x"d6",x"e2",x"c2"),
   469 => (x"87",x"c9",x"c0",x"02"),
   470 => (x"30",x"c4",x"48",x"74"),
   471 => (x"c9",x"c0",x"7e",x"70"),
   472 => (x"f3",x"e6",x"c2",x"87"),
   473 => (x"30",x"c4",x"48",x"bf"),
   474 => (x"e2",x"c2",x"7e",x"70"),
   475 => (x"78",x"6e",x"48",x"da"),
   476 => (x"8e",x"f8",x"48",x"c1"),
   477 => (x"4c",x"26",x"4d",x"26"),
   478 => (x"4f",x"26",x"4b",x"26"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"4a",x"71",x"0e",x"5d"),
   481 => (x"bf",x"d6",x"e2",x"c2"),
   482 => (x"72",x"87",x"cb",x"02"),
   483 => (x"72",x"2b",x"c7",x"4b"),
   484 => (x"9c",x"ff",x"c1",x"4c"),
   485 => (x"4b",x"72",x"87",x"c9"),
   486 => (x"4c",x"72",x"2b",x"c8"),
   487 => (x"c2",x"9c",x"ff",x"c3"),
   488 => (x"83",x"bf",x"e3",x"e6"),
   489 => (x"bf",x"dc",x"f0",x"c0"),
   490 => (x"87",x"d9",x"02",x"ab"),
   491 => (x"5b",x"e0",x"f0",x"c0"),
   492 => (x"1e",x"ce",x"da",x"c2"),
   493 => (x"fd",x"f0",x"49",x"73"),
   494 => (x"70",x"86",x"c4",x"87"),
   495 => (x"87",x"c5",x"05",x"98"),
   496 => (x"e6",x"c0",x"48",x"c0"),
   497 => (x"d6",x"e2",x"c2",x"87"),
   498 => (x"87",x"d2",x"02",x"bf"),
   499 => (x"91",x"c4",x"49",x"74"),
   500 => (x"81",x"ce",x"da",x"c2"),
   501 => (x"ff",x"cf",x"4d",x"69"),
   502 => (x"9d",x"ff",x"ff",x"ff"),
   503 => (x"49",x"74",x"87",x"cb"),
   504 => (x"da",x"c2",x"91",x"c2"),
   505 => (x"69",x"9f",x"81",x"ce"),
   506 => (x"fe",x"48",x"75",x"4d"),
   507 => (x"5e",x"0e",x"87",x"c6"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"c0",x"4d",x"71",x"1e"),
   510 => (x"c9",x"49",x"c1",x"1e"),
   511 => (x"86",x"c4",x"87",x"c7"),
   512 => (x"02",x"9c",x"4c",x"70"),
   513 => (x"c2",x"87",x"c0",x"c1"),
   514 => (x"75",x"4a",x"de",x"e2"),
   515 => (x"87",x"ff",x"e0",x"49"),
   516 => (x"c0",x"02",x"98",x"70"),
   517 => (x"4a",x"74",x"87",x"f1"),
   518 => (x"4b",x"cb",x"49",x"75"),
   519 => (x"70",x"87",x"e5",x"e1"),
   520 => (x"e2",x"c0",x"02",x"98"),
   521 => (x"74",x"1e",x"c0",x"87"),
   522 => (x"87",x"c7",x"02",x"9c"),
   523 => (x"c0",x"48",x"a6",x"c4"),
   524 => (x"c4",x"87",x"c5",x"78"),
   525 => (x"78",x"c1",x"48",x"a6"),
   526 => (x"c8",x"49",x"66",x"c4"),
   527 => (x"86",x"c4",x"87",x"c7"),
   528 => (x"05",x"9c",x"4c",x"70"),
   529 => (x"74",x"87",x"c0",x"ff"),
   530 => (x"e7",x"fc",x"26",x"48"),
   531 => (x"5b",x"5e",x"0e",x"87"),
   532 => (x"1e",x"0e",x"5d",x"5c"),
   533 => (x"05",x"9b",x"4b",x"71"),
   534 => (x"48",x"c0",x"87",x"c5"),
   535 => (x"c8",x"87",x"e5",x"c1"),
   536 => (x"7d",x"c0",x"4d",x"a3"),
   537 => (x"c7",x"02",x"66",x"d4"),
   538 => (x"97",x"66",x"d4",x"87"),
   539 => (x"87",x"c5",x"05",x"bf"),
   540 => (x"cf",x"c1",x"48",x"c0"),
   541 => (x"49",x"66",x"d4",x"87"),
   542 => (x"70",x"87",x"f3",x"fd"),
   543 => (x"c1",x"02",x"9c",x"4c"),
   544 => (x"a4",x"dc",x"87",x"c0"),
   545 => (x"da",x"7d",x"69",x"49"),
   546 => (x"a3",x"c4",x"49",x"a4"),
   547 => (x"7a",x"69",x"9f",x"4a"),
   548 => (x"bf",x"d6",x"e2",x"c2"),
   549 => (x"d4",x"87",x"d2",x"02"),
   550 => (x"69",x"9f",x"49",x"a4"),
   551 => (x"ff",x"ff",x"c0",x"49"),
   552 => (x"d0",x"48",x"71",x"99"),
   553 => (x"c2",x"7e",x"70",x"30"),
   554 => (x"6e",x"7e",x"c0",x"87"),
   555 => (x"80",x"6a",x"48",x"49"),
   556 => (x"7b",x"c0",x"7a",x"70"),
   557 => (x"6a",x"49",x"a3",x"cc"),
   558 => (x"49",x"a3",x"d0",x"79"),
   559 => (x"48",x"74",x"79",x"c0"),
   560 => (x"48",x"c0",x"87",x"c2"),
   561 => (x"87",x"ec",x"fa",x"26"),
   562 => (x"5c",x"5b",x"5e",x"0e"),
   563 => (x"4c",x"71",x"0e",x"5d"),
   564 => (x"48",x"dc",x"f0",x"c0"),
   565 => (x"9c",x"74",x"78",x"ff"),
   566 => (x"87",x"ca",x"c1",x"02"),
   567 => (x"69",x"49",x"a4",x"c8"),
   568 => (x"87",x"c2",x"c1",x"02"),
   569 => (x"6c",x"4a",x"66",x"d0"),
   570 => (x"a6",x"d4",x"82",x"49"),
   571 => (x"4d",x"66",x"d0",x"5a"),
   572 => (x"d2",x"e2",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e4",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"f4",x"f9",x"49"),
   578 => (x"e2",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"ce"),
   580 => (x"75",x"7c",x"71",x"81"),
   581 => (x"d2",x"e2",x"c2",x"b9"),
   582 => (x"ba",x"ff",x"4a",x"bf"),
   583 => (x"99",x"71",x"99",x"72"),
   584 => (x"87",x"dc",x"ff",x"05"),
   585 => (x"cb",x"f9",x"7c",x"75"),
   586 => (x"1e",x"73",x"1e",x"87"),
   587 => (x"02",x"9b",x"4b",x"71"),
   588 => (x"a3",x"c8",x"87",x"c7"),
   589 => (x"c5",x"05",x"69",x"49"),
   590 => (x"c0",x"48",x"c0",x"87"),
   591 => (x"e6",x"c2",x"87",x"eb"),
   592 => (x"c4",x"4a",x"bf",x"e7"),
   593 => (x"49",x"69",x"49",x"a3"),
   594 => (x"e2",x"c2",x"89",x"c2"),
   595 => (x"71",x"91",x"bf",x"ce"),
   596 => (x"e2",x"c2",x"4a",x"a2"),
   597 => (x"6b",x"49",x"bf",x"d2"),
   598 => (x"4a",x"a2",x"71",x"99"),
   599 => (x"72",x"1e",x"66",x"c8"),
   600 => (x"87",x"d2",x"ea",x"49"),
   601 => (x"49",x"70",x"86",x"c4"),
   602 => (x"87",x"cc",x"f8",x"48"),
   603 => (x"71",x"1e",x"73",x"1e"),
   604 => (x"c7",x"02",x"9b",x"4b"),
   605 => (x"49",x"a3",x"c8",x"87"),
   606 => (x"87",x"c5",x"05",x"69"),
   607 => (x"eb",x"c0",x"48",x"c0"),
   608 => (x"e7",x"e6",x"c2",x"87"),
   609 => (x"a3",x"c4",x"4a",x"bf"),
   610 => (x"c2",x"49",x"69",x"49"),
   611 => (x"ce",x"e2",x"c2",x"89"),
   612 => (x"a2",x"71",x"91",x"bf"),
   613 => (x"d2",x"e2",x"c2",x"4a"),
   614 => (x"99",x"6b",x"49",x"bf"),
   615 => (x"c8",x"4a",x"a2",x"71"),
   616 => (x"49",x"72",x"1e",x"66"),
   617 => (x"c4",x"87",x"c5",x"e6"),
   618 => (x"48",x"49",x"70",x"86"),
   619 => (x"1e",x"87",x"c9",x"f7"),
   620 => (x"4b",x"71",x"1e",x"73"),
   621 => (x"e4",x"c0",x"02",x"9b"),
   622 => (x"fb",x"e6",x"c2",x"87"),
   623 => (x"c2",x"4a",x"73",x"5b"),
   624 => (x"ce",x"e2",x"c2",x"8a"),
   625 => (x"c2",x"92",x"49",x"bf"),
   626 => (x"48",x"bf",x"e7",x"e6"),
   627 => (x"e6",x"c2",x"80",x"72"),
   628 => (x"48",x"71",x"58",x"ff"),
   629 => (x"e2",x"c2",x"30",x"c4"),
   630 => (x"ed",x"c0",x"58",x"de"),
   631 => (x"f7",x"e6",x"c2",x"87"),
   632 => (x"eb",x"e6",x"c2",x"48"),
   633 => (x"e6",x"c2",x"78",x"bf"),
   634 => (x"e6",x"c2",x"48",x"fb"),
   635 => (x"c2",x"78",x"bf",x"ef"),
   636 => (x"02",x"bf",x"d6",x"e2"),
   637 => (x"e2",x"c2",x"87",x"c9"),
   638 => (x"c4",x"49",x"bf",x"ce"),
   639 => (x"c2",x"87",x"c7",x"31"),
   640 => (x"49",x"bf",x"f3",x"e6"),
   641 => (x"e2",x"c2",x"31",x"c4"),
   642 => (x"eb",x"f5",x"59",x"de"),
   643 => (x"5b",x"5e",x"0e",x"87"),
   644 => (x"4a",x"71",x"0e",x"5c"),
   645 => (x"9a",x"72",x"4b",x"c0"),
   646 => (x"87",x"e1",x"c0",x"02"),
   647 => (x"9f",x"49",x"a2",x"da"),
   648 => (x"e2",x"c2",x"4b",x"69"),
   649 => (x"cf",x"02",x"bf",x"d6"),
   650 => (x"49",x"a2",x"d4",x"87"),
   651 => (x"4c",x"49",x"69",x"9f"),
   652 => (x"9c",x"ff",x"ff",x"c0"),
   653 => (x"87",x"c2",x"34",x"d0"),
   654 => (x"49",x"74",x"4c",x"c0"),
   655 => (x"fd",x"49",x"73",x"b3"),
   656 => (x"f1",x"f4",x"87",x"ed"),
   657 => (x"5b",x"5e",x"0e",x"87"),
   658 => (x"f4",x"0e",x"5d",x"5c"),
   659 => (x"c0",x"4a",x"71",x"86"),
   660 => (x"02",x"9a",x"72",x"7e"),
   661 => (x"da",x"c2",x"87",x"d8"),
   662 => (x"78",x"c0",x"48",x"ca"),
   663 => (x"48",x"c2",x"da",x"c2"),
   664 => (x"bf",x"fb",x"e6",x"c2"),
   665 => (x"c6",x"da",x"c2",x"78"),
   666 => (x"f7",x"e6",x"c2",x"48"),
   667 => (x"e2",x"c2",x"78",x"bf"),
   668 => (x"50",x"c0",x"48",x"eb"),
   669 => (x"bf",x"da",x"e2",x"c2"),
   670 => (x"ca",x"da",x"c2",x"49"),
   671 => (x"aa",x"71",x"4a",x"bf"),
   672 => (x"87",x"ff",x"c3",x"03"),
   673 => (x"99",x"cf",x"49",x"72"),
   674 => (x"87",x"e0",x"c0",x"05"),
   675 => (x"1e",x"ce",x"da",x"c2"),
   676 => (x"bf",x"c2",x"da",x"c2"),
   677 => (x"c2",x"da",x"c2",x"49"),
   678 => (x"78",x"a1",x"c1",x"48"),
   679 => (x"87",x"d6",x"e5",x"71"),
   680 => (x"f0",x"c0",x"86",x"c4"),
   681 => (x"da",x"c2",x"48",x"d8"),
   682 => (x"87",x"cc",x"78",x"ce"),
   683 => (x"bf",x"d8",x"f0",x"c0"),
   684 => (x"80",x"e0",x"c0",x"48"),
   685 => (x"58",x"dc",x"f0",x"c0"),
   686 => (x"bf",x"ca",x"da",x"c2"),
   687 => (x"c2",x"80",x"c1",x"48"),
   688 => (x"27",x"58",x"ce",x"da"),
   689 => (x"00",x"00",x"0c",x"18"),
   690 => (x"4d",x"bf",x"97",x"bf"),
   691 => (x"e2",x"c2",x"02",x"9d"),
   692 => (x"ad",x"e5",x"c3",x"87"),
   693 => (x"87",x"db",x"c2",x"02"),
   694 => (x"bf",x"d8",x"f0",x"c0"),
   695 => (x"49",x"a3",x"cb",x"4b"),
   696 => (x"ac",x"cf",x"4c",x"11"),
   697 => (x"87",x"d2",x"c1",x"05"),
   698 => (x"99",x"df",x"49",x"75"),
   699 => (x"91",x"cd",x"89",x"c1"),
   700 => (x"81",x"de",x"e2",x"c2"),
   701 => (x"12",x"4a",x"a3",x"c1"),
   702 => (x"4a",x"a3",x"c3",x"51"),
   703 => (x"a3",x"c5",x"51",x"12"),
   704 => (x"c7",x"51",x"12",x"4a"),
   705 => (x"51",x"12",x"4a",x"a3"),
   706 => (x"12",x"4a",x"a3",x"c9"),
   707 => (x"4a",x"a3",x"ce",x"51"),
   708 => (x"a3",x"d0",x"51",x"12"),
   709 => (x"d2",x"51",x"12",x"4a"),
   710 => (x"51",x"12",x"4a",x"a3"),
   711 => (x"12",x"4a",x"a3",x"d4"),
   712 => (x"4a",x"a3",x"d6",x"51"),
   713 => (x"a3",x"d8",x"51",x"12"),
   714 => (x"dc",x"51",x"12",x"4a"),
   715 => (x"51",x"12",x"4a",x"a3"),
   716 => (x"12",x"4a",x"a3",x"de"),
   717 => (x"c0",x"7e",x"c1",x"51"),
   718 => (x"49",x"74",x"87",x"f9"),
   719 => (x"c0",x"05",x"99",x"c8"),
   720 => (x"49",x"74",x"87",x"ea"),
   721 => (x"d0",x"05",x"99",x"d0"),
   722 => (x"02",x"66",x"dc",x"87"),
   723 => (x"73",x"87",x"ca",x"c0"),
   724 => (x"0f",x"66",x"dc",x"49"),
   725 => (x"d3",x"02",x"98",x"70"),
   726 => (x"c0",x"05",x"6e",x"87"),
   727 => (x"e2",x"c2",x"87",x"c6"),
   728 => (x"50",x"c0",x"48",x"de"),
   729 => (x"bf",x"d8",x"f0",x"c0"),
   730 => (x"87",x"e7",x"c2",x"48"),
   731 => (x"48",x"eb",x"e2",x"c2"),
   732 => (x"c2",x"7e",x"50",x"c0"),
   733 => (x"49",x"bf",x"da",x"e2"),
   734 => (x"bf",x"ca",x"da",x"c2"),
   735 => (x"04",x"aa",x"71",x"4a"),
   736 => (x"c2",x"87",x"c1",x"fc"),
   737 => (x"05",x"bf",x"fb",x"e6"),
   738 => (x"c2",x"87",x"c8",x"c0"),
   739 => (x"02",x"bf",x"d6",x"e2"),
   740 => (x"c0",x"87",x"fe",x"c1"),
   741 => (x"ff",x"48",x"dc",x"f0"),
   742 => (x"c6",x"da",x"c2",x"78"),
   743 => (x"db",x"ef",x"49",x"bf"),
   744 => (x"c2",x"49",x"70",x"87"),
   745 => (x"c4",x"59",x"ca",x"da"),
   746 => (x"da",x"c2",x"48",x"a6"),
   747 => (x"c2",x"78",x"bf",x"c6"),
   748 => (x"02",x"bf",x"d6",x"e2"),
   749 => (x"c4",x"87",x"d8",x"c0"),
   750 => (x"ff",x"cf",x"49",x"66"),
   751 => (x"99",x"f8",x"ff",x"ff"),
   752 => (x"c5",x"c0",x"02",x"a9"),
   753 => (x"c0",x"4d",x"c0",x"87"),
   754 => (x"4d",x"c1",x"87",x"e1"),
   755 => (x"c4",x"87",x"dc",x"c0"),
   756 => (x"ff",x"cf",x"49",x"66"),
   757 => (x"02",x"a9",x"99",x"f8"),
   758 => (x"c8",x"87",x"c8",x"c0"),
   759 => (x"78",x"c0",x"48",x"a6"),
   760 => (x"c8",x"87",x"c5",x"c0"),
   761 => (x"78",x"c1",x"48",x"a6"),
   762 => (x"75",x"4d",x"66",x"c8"),
   763 => (x"e0",x"c0",x"05",x"9d"),
   764 => (x"49",x"66",x"c4",x"87"),
   765 => (x"e2",x"c2",x"89",x"c2"),
   766 => (x"91",x"4a",x"bf",x"ce"),
   767 => (x"bf",x"e7",x"e6",x"c2"),
   768 => (x"c2",x"da",x"c2",x"4a"),
   769 => (x"78",x"a1",x"72",x"48"),
   770 => (x"48",x"ca",x"da",x"c2"),
   771 => (x"e3",x"f9",x"78",x"c0"),
   772 => (x"f4",x"48",x"c0",x"87"),
   773 => (x"87",x"dc",x"ed",x"8e"),
   774 => (x"00",x"00",x"00",x"00"),
   775 => (x"ff",x"ff",x"ff",x"ff"),
   776 => (x"00",x"00",x"0c",x"28"),
   777 => (x"00",x"00",x"0c",x"31"),
   778 => (x"33",x"54",x"41",x"46"),
   779 => (x"20",x"20",x"20",x"32"),
   780 => (x"54",x"41",x"46",x"00"),
   781 => (x"20",x"20",x"36",x"31"),
   782 => (x"ff",x"1e",x"00",x"20"),
   783 => (x"ff",x"c3",x"48",x"d4"),
   784 => (x"26",x"48",x"68",x"78"),
   785 => (x"d4",x"ff",x"1e",x"4f"),
   786 => (x"78",x"ff",x"c3",x"48"),
   787 => (x"c8",x"48",x"d0",x"ff"),
   788 => (x"d4",x"ff",x"78",x"e1"),
   789 => (x"c2",x"78",x"d4",x"48"),
   790 => (x"ff",x"48",x"ff",x"e6"),
   791 => (x"26",x"50",x"bf",x"d4"),
   792 => (x"d0",x"ff",x"1e",x"4f"),
   793 => (x"78",x"e0",x"c0",x"48"),
   794 => (x"ff",x"1e",x"4f",x"26"),
   795 => (x"49",x"70",x"87",x"cc"),
   796 => (x"87",x"c6",x"02",x"99"),
   797 => (x"05",x"a9",x"fb",x"c0"),
   798 => (x"48",x"71",x"87",x"f1"),
   799 => (x"5e",x"0e",x"4f",x"26"),
   800 => (x"71",x"0e",x"5c",x"5b"),
   801 => (x"fe",x"4c",x"c0",x"4b"),
   802 => (x"49",x"70",x"87",x"f0"),
   803 => (x"f9",x"c0",x"02",x"99"),
   804 => (x"a9",x"ec",x"c0",x"87"),
   805 => (x"87",x"f2",x"c0",x"02"),
   806 => (x"02",x"a9",x"fb",x"c0"),
   807 => (x"cc",x"87",x"eb",x"c0"),
   808 => (x"03",x"ac",x"b7",x"66"),
   809 => (x"66",x"d0",x"87",x"c7"),
   810 => (x"71",x"87",x"c2",x"02"),
   811 => (x"02",x"99",x"71",x"53"),
   812 => (x"84",x"c1",x"87",x"c2"),
   813 => (x"70",x"87",x"c3",x"fe"),
   814 => (x"cd",x"02",x"99",x"49"),
   815 => (x"a9",x"ec",x"c0",x"87"),
   816 => (x"c0",x"87",x"c7",x"02"),
   817 => (x"ff",x"05",x"a9",x"fb"),
   818 => (x"66",x"d0",x"87",x"d5"),
   819 => (x"c0",x"87",x"c3",x"02"),
   820 => (x"ec",x"c0",x"7b",x"97"),
   821 => (x"87",x"c4",x"05",x"a9"),
   822 => (x"87",x"c5",x"4a",x"74"),
   823 => (x"0a",x"c0",x"4a",x"74"),
   824 => (x"c2",x"48",x"72",x"8a"),
   825 => (x"26",x"4d",x"26",x"87"),
   826 => (x"26",x"4b",x"26",x"4c"),
   827 => (x"c9",x"fd",x"1e",x"4f"),
   828 => (x"c0",x"49",x"70",x"87"),
   829 => (x"04",x"a9",x"b7",x"f0"),
   830 => (x"f9",x"c0",x"87",x"ca"),
   831 => (x"c3",x"01",x"a9",x"b7"),
   832 => (x"89",x"f0",x"c0",x"87"),
   833 => (x"a9",x"b7",x"c1",x"c1"),
   834 => (x"c1",x"87",x"ca",x"04"),
   835 => (x"01",x"a9",x"b7",x"da"),
   836 => (x"f7",x"c0",x"87",x"c3"),
   837 => (x"26",x"48",x"71",x"89"),
   838 => (x"5b",x"5e",x"0e",x"4f"),
   839 => (x"4a",x"71",x"0e",x"5c"),
   840 => (x"72",x"4c",x"d4",x"ff"),
   841 => (x"87",x"ea",x"c0",x"49"),
   842 => (x"02",x"9b",x"4b",x"70"),
   843 => (x"8b",x"c1",x"87",x"c2"),
   844 => (x"c8",x"48",x"d0",x"ff"),
   845 => (x"d5",x"c1",x"78",x"c5"),
   846 => (x"c6",x"49",x"73",x"7c"),
   847 => (x"fa",x"d5",x"c2",x"31"),
   848 => (x"48",x"4a",x"bf",x"97"),
   849 => (x"7c",x"70",x"b0",x"71"),
   850 => (x"c4",x"48",x"d0",x"ff"),
   851 => (x"fe",x"48",x"73",x"78"),
   852 => (x"5e",x"0e",x"87",x"d5"),
   853 => (x"0e",x"5d",x"5c",x"5b"),
   854 => (x"4b",x"71",x"86",x"f8"),
   855 => (x"f8",x"c0",x"7e",x"c0"),
   856 => (x"49",x"bf",x"97",x"f9"),
   857 => (x"c0",x"05",x"a9",x"df"),
   858 => (x"a3",x"c8",x"87",x"ee"),
   859 => (x"49",x"69",x"97",x"49"),
   860 => (x"05",x"a9",x"c3",x"c1"),
   861 => (x"a3",x"c9",x"87",x"dd"),
   862 => (x"49",x"69",x"97",x"49"),
   863 => (x"05",x"a9",x"c6",x"c1"),
   864 => (x"a3",x"ca",x"87",x"d1"),
   865 => (x"49",x"69",x"97",x"49"),
   866 => (x"05",x"a9",x"c7",x"c1"),
   867 => (x"48",x"c1",x"87",x"c5"),
   868 => (x"c0",x"87",x"e1",x"c2"),
   869 => (x"87",x"dc",x"c2",x"48"),
   870 => (x"c0",x"87",x"ea",x"fa"),
   871 => (x"f9",x"f8",x"c0",x"4c"),
   872 => (x"c0",x"49",x"bf",x"97"),
   873 => (x"87",x"cf",x"04",x"a9"),
   874 => (x"c1",x"87",x"ff",x"fa"),
   875 => (x"f9",x"f8",x"c0",x"84"),
   876 => (x"ac",x"49",x"bf",x"97"),
   877 => (x"c0",x"87",x"f1",x"06"),
   878 => (x"bf",x"97",x"f9",x"f8"),
   879 => (x"f9",x"87",x"cf",x"02"),
   880 => (x"49",x"70",x"87",x"f8"),
   881 => (x"87",x"c6",x"02",x"99"),
   882 => (x"05",x"a9",x"ec",x"c0"),
   883 => (x"4c",x"c0",x"87",x"f1"),
   884 => (x"70",x"87",x"e7",x"f9"),
   885 => (x"87",x"e2",x"f9",x"4d"),
   886 => (x"f9",x"58",x"a6",x"c8"),
   887 => (x"4a",x"70",x"87",x"dc"),
   888 => (x"a3",x"c8",x"84",x"c1"),
   889 => (x"49",x"69",x"97",x"49"),
   890 => (x"87",x"c7",x"02",x"ad"),
   891 => (x"05",x"ad",x"ff",x"c0"),
   892 => (x"c9",x"87",x"e7",x"c0"),
   893 => (x"69",x"97",x"49",x"a3"),
   894 => (x"a9",x"66",x"c4",x"49"),
   895 => (x"48",x"87",x"c7",x"02"),
   896 => (x"05",x"a8",x"ff",x"c0"),
   897 => (x"a3",x"ca",x"87",x"d4"),
   898 => (x"49",x"69",x"97",x"49"),
   899 => (x"87",x"c6",x"02",x"aa"),
   900 => (x"05",x"aa",x"ff",x"c0"),
   901 => (x"7e",x"c1",x"87",x"c4"),
   902 => (x"ec",x"c0",x"87",x"d0"),
   903 => (x"87",x"c6",x"02",x"ad"),
   904 => (x"05",x"ad",x"fb",x"c0"),
   905 => (x"4c",x"c0",x"87",x"c4"),
   906 => (x"02",x"6e",x"7e",x"c1"),
   907 => (x"f8",x"87",x"e1",x"fe"),
   908 => (x"48",x"74",x"87",x"ef"),
   909 => (x"ec",x"fa",x"8e",x"f8"),
   910 => (x"5e",x"0e",x"00",x"87"),
   911 => (x"0e",x"5d",x"5c",x"5b"),
   912 => (x"c0",x"4b",x"71",x"1e"),
   913 => (x"04",x"ab",x"4d",x"4c"),
   914 => (x"c0",x"87",x"e8",x"c0"),
   915 => (x"75",x"1e",x"d2",x"f5"),
   916 => (x"87",x"c4",x"02",x"9d"),
   917 => (x"87",x"c2",x"4a",x"c0"),
   918 => (x"49",x"72",x"4a",x"c1"),
   919 => (x"c4",x"87",x"e6",x"ef"),
   920 => (x"c1",x"7e",x"70",x"86"),
   921 => (x"c2",x"05",x"6e",x"84"),
   922 => (x"c1",x"4c",x"73",x"87"),
   923 => (x"06",x"ac",x"73",x"85"),
   924 => (x"6e",x"87",x"d8",x"ff"),
   925 => (x"4d",x"26",x"26",x"48"),
   926 => (x"4b",x"26",x"4c",x"26"),
   927 => (x"5e",x"0e",x"4f",x"26"),
   928 => (x"0e",x"5d",x"5c",x"5b"),
   929 => (x"49",x"4c",x"71",x"1e"),
   930 => (x"e7",x"c2",x"91",x"de"),
   931 => (x"85",x"71",x"4d",x"d9"),
   932 => (x"c1",x"02",x"6d",x"97"),
   933 => (x"e7",x"c2",x"87",x"dd"),
   934 => (x"74",x"4a",x"bf",x"c4"),
   935 => (x"fe",x"49",x"72",x"82"),
   936 => (x"7e",x"70",x"87",x"d8"),
   937 => (x"f3",x"c0",x"02",x"6e"),
   938 => (x"cc",x"e7",x"c2",x"87"),
   939 => (x"cb",x"4a",x"6e",x"4b"),
   940 => (x"f3",x"c7",x"ff",x"49"),
   941 => (x"cb",x"4b",x"74",x"87"),
   942 => (x"f2",x"e0",x"c1",x"93"),
   943 => (x"c0",x"83",x"c4",x"83"),
   944 => (x"74",x"7b",x"f7",x"fb"),
   945 => (x"f4",x"c6",x"c1",x"49"),
   946 => (x"c2",x"7b",x"75",x"87"),
   947 => (x"bf",x"97",x"d8",x"e7"),
   948 => (x"e7",x"c2",x"1e",x"49"),
   949 => (x"d9",x"c1",x"49",x"cc"),
   950 => (x"86",x"c4",x"87",x"f2"),
   951 => (x"c6",x"c1",x"49",x"74"),
   952 => (x"49",x"c0",x"87",x"db"),
   953 => (x"87",x"fa",x"c7",x"c1"),
   954 => (x"48",x"c0",x"e7",x"c2"),
   955 => (x"49",x"c1",x"78",x"c0"),
   956 => (x"26",x"87",x"fd",x"df"),
   957 => (x"4c",x"87",x"ff",x"fd"),
   958 => (x"69",x"64",x"61",x"6f"),
   959 => (x"2e",x"2e",x"67",x"6e"),
   960 => (x"5e",x"0e",x"00",x"2e"),
   961 => (x"71",x"0e",x"5c",x"5b"),
   962 => (x"e7",x"c2",x"4a",x"4b"),
   963 => (x"72",x"82",x"bf",x"c4"),
   964 => (x"87",x"e6",x"fc",x"49"),
   965 => (x"02",x"9c",x"4c",x"70"),
   966 => (x"eb",x"49",x"87",x"c4"),
   967 => (x"e7",x"c2",x"87",x"ef"),
   968 => (x"78",x"c0",x"48",x"c4"),
   969 => (x"c7",x"df",x"49",x"c1"),
   970 => (x"87",x"cc",x"fd",x"87"),
   971 => (x"5c",x"5b",x"5e",x"0e"),
   972 => (x"86",x"f4",x"0e",x"5d"),
   973 => (x"4d",x"ce",x"da",x"c2"),
   974 => (x"a6",x"c4",x"4c",x"c0"),
   975 => (x"c2",x"78",x"c0",x"48"),
   976 => (x"49",x"bf",x"c4",x"e7"),
   977 => (x"c1",x"06",x"a9",x"c0"),
   978 => (x"da",x"c2",x"87",x"c1"),
   979 => (x"02",x"98",x"48",x"ce"),
   980 => (x"c0",x"87",x"f8",x"c0"),
   981 => (x"c8",x"1e",x"d2",x"f5"),
   982 => (x"87",x"c7",x"02",x"66"),
   983 => (x"c0",x"48",x"a6",x"c4"),
   984 => (x"c4",x"87",x"c5",x"78"),
   985 => (x"78",x"c1",x"48",x"a6"),
   986 => (x"eb",x"49",x"66",x"c4"),
   987 => (x"86",x"c4",x"87",x"d7"),
   988 => (x"84",x"c1",x"4d",x"70"),
   989 => (x"c1",x"48",x"66",x"c4"),
   990 => (x"58",x"a6",x"c8",x"80"),
   991 => (x"bf",x"c4",x"e7",x"c2"),
   992 => (x"c6",x"03",x"ac",x"49"),
   993 => (x"05",x"9d",x"75",x"87"),
   994 => (x"c0",x"87",x"c8",x"ff"),
   995 => (x"02",x"9d",x"75",x"4c"),
   996 => (x"c0",x"87",x"e0",x"c3"),
   997 => (x"c8",x"1e",x"d2",x"f5"),
   998 => (x"87",x"c7",x"02",x"66"),
   999 => (x"c0",x"48",x"a6",x"cc"),
  1000 => (x"cc",x"87",x"c5",x"78"),
  1001 => (x"78",x"c1",x"48",x"a6"),
  1002 => (x"ea",x"49",x"66",x"cc"),
  1003 => (x"86",x"c4",x"87",x"d7"),
  1004 => (x"02",x"6e",x"7e",x"70"),
  1005 => (x"6e",x"87",x"e9",x"c2"),
  1006 => (x"97",x"81",x"cb",x"49"),
  1007 => (x"99",x"d0",x"49",x"69"),
  1008 => (x"87",x"d6",x"c1",x"02"),
  1009 => (x"4a",x"c2",x"fc",x"c0"),
  1010 => (x"91",x"cb",x"49",x"74"),
  1011 => (x"81",x"f2",x"e0",x"c1"),
  1012 => (x"81",x"c8",x"79",x"72"),
  1013 => (x"74",x"51",x"ff",x"c3"),
  1014 => (x"c2",x"91",x"de",x"49"),
  1015 => (x"71",x"4d",x"d9",x"e7"),
  1016 => (x"97",x"c1",x"c2",x"85"),
  1017 => (x"49",x"a5",x"c1",x"7d"),
  1018 => (x"c2",x"51",x"e0",x"c0"),
  1019 => (x"bf",x"97",x"de",x"e2"),
  1020 => (x"c1",x"87",x"d2",x"02"),
  1021 => (x"4b",x"a5",x"c2",x"84"),
  1022 => (x"4a",x"de",x"e2",x"c2"),
  1023 => (x"c2",x"ff",x"49",x"db"),
  1024 => (x"db",x"c1",x"87",x"e6"),
  1025 => (x"49",x"a5",x"cd",x"87"),
  1026 => (x"84",x"c1",x"51",x"c0"),
  1027 => (x"6e",x"4b",x"a5",x"c2"),
  1028 => (x"ff",x"49",x"cb",x"4a"),
  1029 => (x"c1",x"87",x"d1",x"c2"),
  1030 => (x"f9",x"c0",x"87",x"c6"),
  1031 => (x"49",x"74",x"4a",x"fe"),
  1032 => (x"e0",x"c1",x"91",x"cb"),
  1033 => (x"79",x"72",x"81",x"f2"),
  1034 => (x"97",x"de",x"e2",x"c2"),
  1035 => (x"87",x"d8",x"02",x"bf"),
  1036 => (x"91",x"de",x"49",x"74"),
  1037 => (x"e7",x"c2",x"84",x"c1"),
  1038 => (x"83",x"71",x"4b",x"d9"),
  1039 => (x"4a",x"de",x"e2",x"c2"),
  1040 => (x"c1",x"ff",x"49",x"dd"),
  1041 => (x"87",x"d8",x"87",x"e2"),
  1042 => (x"93",x"de",x"4b",x"74"),
  1043 => (x"83",x"d9",x"e7",x"c2"),
  1044 => (x"c0",x"49",x"a3",x"cb"),
  1045 => (x"73",x"84",x"c1",x"51"),
  1046 => (x"49",x"cb",x"4a",x"6e"),
  1047 => (x"87",x"c8",x"c1",x"ff"),
  1048 => (x"c1",x"48",x"66",x"c4"),
  1049 => (x"58",x"a6",x"c8",x"80"),
  1050 => (x"c0",x"03",x"ac",x"c7"),
  1051 => (x"05",x"6e",x"87",x"c5"),
  1052 => (x"74",x"87",x"e0",x"fc"),
  1053 => (x"f7",x"8e",x"f4",x"48"),
  1054 => (x"73",x"1e",x"87",x"fc"),
  1055 => (x"49",x"4b",x"71",x"1e"),
  1056 => (x"e0",x"c1",x"91",x"cb"),
  1057 => (x"a1",x"c8",x"81",x"f2"),
  1058 => (x"fa",x"d5",x"c2",x"4a"),
  1059 => (x"c9",x"50",x"12",x"48"),
  1060 => (x"f8",x"c0",x"4a",x"a1"),
  1061 => (x"50",x"12",x"48",x"f9"),
  1062 => (x"e7",x"c2",x"81",x"ca"),
  1063 => (x"50",x"11",x"48",x"d8"),
  1064 => (x"97",x"d8",x"e7",x"c2"),
  1065 => (x"c0",x"1e",x"49",x"bf"),
  1066 => (x"df",x"d2",x"c1",x"49"),
  1067 => (x"c0",x"e7",x"c2",x"87"),
  1068 => (x"c1",x"78",x"de",x"48"),
  1069 => (x"87",x"f8",x"d8",x"49"),
  1070 => (x"87",x"fe",x"f6",x"26"),
  1071 => (x"49",x"4a",x"71",x"1e"),
  1072 => (x"e0",x"c1",x"91",x"cb"),
  1073 => (x"81",x"c8",x"81",x"f2"),
  1074 => (x"e7",x"c2",x"48",x"11"),
  1075 => (x"e7",x"c2",x"58",x"c4"),
  1076 => (x"78",x"c0",x"48",x"c4"),
  1077 => (x"d7",x"d8",x"49",x"c1"),
  1078 => (x"1e",x"4f",x"26",x"87"),
  1079 => (x"c0",x"c1",x"49",x"c0"),
  1080 => (x"4f",x"26",x"87",x"c0"),
  1081 => (x"02",x"99",x"71",x"1e"),
  1082 => (x"e2",x"c1",x"87",x"d2"),
  1083 => (x"50",x"c0",x"48",x"c7"),
  1084 => (x"c2",x"c1",x"80",x"f7"),
  1085 => (x"e0",x"c1",x"40",x"fc"),
  1086 => (x"87",x"ce",x"78",x"e0"),
  1087 => (x"48",x"c3",x"e2",x"c1"),
  1088 => (x"78",x"c1",x"e0",x"c1"),
  1089 => (x"c3",x"c1",x"80",x"fc"),
  1090 => (x"4f",x"26",x"78",x"db"),
  1091 => (x"5c",x"5b",x"5e",x"0e"),
  1092 => (x"4a",x"4c",x"71",x"0e"),
  1093 => (x"e0",x"c1",x"92",x"cb"),
  1094 => (x"a2",x"c8",x"82",x"f2"),
  1095 => (x"4b",x"a2",x"c9",x"49"),
  1096 => (x"1e",x"4b",x"6b",x"97"),
  1097 => (x"1e",x"49",x"69",x"97"),
  1098 => (x"49",x"12",x"82",x"ca"),
  1099 => (x"87",x"fb",x"ea",x"c0"),
  1100 => (x"fb",x"d6",x"49",x"c0"),
  1101 => (x"c0",x"49",x"74",x"87"),
  1102 => (x"f8",x"87",x"c2",x"fd"),
  1103 => (x"87",x"f8",x"f4",x"8e"),
  1104 => (x"71",x"1e",x"73",x"1e"),
  1105 => (x"c3",x"ff",x"49",x"4b"),
  1106 => (x"fe",x"49",x"73",x"87"),
  1107 => (x"e9",x"f4",x"87",x"fe"),
  1108 => (x"1e",x"73",x"1e",x"87"),
  1109 => (x"a3",x"c6",x"4b",x"71"),
  1110 => (x"87",x"dc",x"02",x"4a"),
  1111 => (x"c0",x"02",x"8a",x"c1"),
  1112 => (x"02",x"8a",x"87",x"e4"),
  1113 => (x"8a",x"87",x"e8",x"c1"),
  1114 => (x"87",x"ca",x"c1",x"02"),
  1115 => (x"ef",x"c0",x"02",x"8a"),
  1116 => (x"d9",x"02",x"8a",x"87"),
  1117 => (x"87",x"e9",x"c1",x"87"),
  1118 => (x"48",x"c0",x"e7",x"c2"),
  1119 => (x"49",x"c1",x"78",x"df"),
  1120 => (x"c1",x"87",x"ed",x"d5"),
  1121 => (x"49",x"c7",x"87",x"e6"),
  1122 => (x"c1",x"87",x"f1",x"fc"),
  1123 => (x"e7",x"c2",x"87",x"de"),
  1124 => (x"c1",x"02",x"bf",x"c4"),
  1125 => (x"c1",x"48",x"87",x"cb"),
  1126 => (x"c8",x"e7",x"c2",x"88"),
  1127 => (x"87",x"c1",x"c1",x"58"),
  1128 => (x"bf",x"c8",x"e7",x"c2"),
  1129 => (x"87",x"f9",x"c0",x"02"),
  1130 => (x"bf",x"c4",x"e7",x"c2"),
  1131 => (x"c2",x"80",x"c1",x"48"),
  1132 => (x"c0",x"58",x"c8",x"e7"),
  1133 => (x"e7",x"c2",x"87",x"eb"),
  1134 => (x"c6",x"49",x"bf",x"c4"),
  1135 => (x"c8",x"e7",x"c2",x"89"),
  1136 => (x"a9",x"b7",x"c0",x"59"),
  1137 => (x"c2",x"87",x"da",x"03"),
  1138 => (x"c0",x"48",x"c4",x"e7"),
  1139 => (x"c2",x"87",x"d2",x"78"),
  1140 => (x"02",x"bf",x"c8",x"e7"),
  1141 => (x"e7",x"c2",x"87",x"cb"),
  1142 => (x"c6",x"48",x"bf",x"c4"),
  1143 => (x"c8",x"e7",x"c2",x"80"),
  1144 => (x"d4",x"49",x"c0",x"58"),
  1145 => (x"49",x"73",x"87",x"ca"),
  1146 => (x"87",x"d1",x"fa",x"c0"),
  1147 => (x"0e",x"87",x"cb",x"f2"),
  1148 => (x"0e",x"5c",x"5b",x"5e"),
  1149 => (x"66",x"cc",x"4c",x"71"),
  1150 => (x"cb",x"4b",x"74",x"1e"),
  1151 => (x"f2",x"e0",x"c1",x"93"),
  1152 => (x"4a",x"a3",x"c4",x"83"),
  1153 => (x"fa",x"fe",x"49",x"6a"),
  1154 => (x"c1",x"c1",x"87",x"ee"),
  1155 => (x"a3",x"c8",x"7b",x"fa"),
  1156 => (x"51",x"66",x"d4",x"49"),
  1157 => (x"d8",x"49",x"a3",x"c9"),
  1158 => (x"a3",x"ca",x"51",x"66"),
  1159 => (x"51",x"66",x"dc",x"49"),
  1160 => (x"87",x"d4",x"f1",x"26"),
  1161 => (x"5c",x"5b",x"5e",x"0e"),
  1162 => (x"d0",x"ff",x"0e",x"5d"),
  1163 => (x"59",x"a6",x"d8",x"86"),
  1164 => (x"c0",x"48",x"a6",x"c8"),
  1165 => (x"c1",x"80",x"fc",x"78"),
  1166 => (x"c8",x"78",x"66",x"c4"),
  1167 => (x"c4",x"78",x"c1",x"80"),
  1168 => (x"c2",x"78",x"c1",x"80"),
  1169 => (x"c1",x"48",x"c8",x"e7"),
  1170 => (x"c0",x"e7",x"c2",x"78"),
  1171 => (x"48",x"6e",x"7e",x"bf"),
  1172 => (x"cb",x"05",x"a8",x"de"),
  1173 => (x"87",x"d4",x"f3",x"87"),
  1174 => (x"a6",x"cc",x"49",x"70"),
  1175 => (x"87",x"f8",x"d0",x"59"),
  1176 => (x"a8",x"df",x"48",x"6e"),
  1177 => (x"87",x"ee",x"c1",x"05"),
  1178 => (x"49",x"66",x"c0",x"c1"),
  1179 => (x"7e",x"69",x"81",x"c4"),
  1180 => (x"48",x"cd",x"db",x"c1"),
  1181 => (x"a1",x"d0",x"49",x"6e"),
  1182 => (x"71",x"41",x"20",x"4a"),
  1183 => (x"87",x"f9",x"05",x"aa"),
  1184 => (x"4a",x"fa",x"c1",x"c1"),
  1185 => (x"0a",x"66",x"c0",x"c1"),
  1186 => (x"c0",x"c1",x"0a",x"7a"),
  1187 => (x"81",x"c9",x"49",x"66"),
  1188 => (x"c0",x"c1",x"51",x"df"),
  1189 => (x"81",x"ca",x"49",x"66"),
  1190 => (x"c1",x"51",x"d3",x"c1"),
  1191 => (x"cb",x"49",x"66",x"c0"),
  1192 => (x"4b",x"a1",x"c4",x"81"),
  1193 => (x"6b",x"48",x"a6",x"c4"),
  1194 => (x"72",x"1e",x"71",x"78"),
  1195 => (x"dd",x"db",x"c1",x"1e"),
  1196 => (x"49",x"66",x"cc",x"48"),
  1197 => (x"20",x"4a",x"a1",x"d0"),
  1198 => (x"05",x"aa",x"71",x"41"),
  1199 => (x"4a",x"26",x"87",x"f9"),
  1200 => (x"79",x"72",x"49",x"26"),
  1201 => (x"df",x"4a",x"a1",x"c9"),
  1202 => (x"c1",x"81",x"ca",x"52"),
  1203 => (x"a6",x"c8",x"51",x"d4"),
  1204 => (x"cf",x"78",x"c2",x"48"),
  1205 => (x"ec",x"e5",x"87",x"c2"),
  1206 => (x"87",x"ce",x"e6",x"87"),
  1207 => (x"70",x"87",x"db",x"e5"),
  1208 => (x"ac",x"fb",x"c0",x"4c"),
  1209 => (x"87",x"d0",x"c1",x"02"),
  1210 => (x"c1",x"05",x"66",x"d4"),
  1211 => (x"1e",x"c0",x"87",x"c2"),
  1212 => (x"c1",x"1e",x"c1",x"1e"),
  1213 => (x"c0",x"1e",x"e5",x"e2"),
  1214 => (x"87",x"f3",x"fb",x"49"),
  1215 => (x"4a",x"66",x"d0",x"c1"),
  1216 => (x"49",x"6a",x"82",x"c4"),
  1217 => (x"51",x"74",x"81",x"c7"),
  1218 => (x"1e",x"d8",x"1e",x"c1"),
  1219 => (x"81",x"c8",x"49",x"6a"),
  1220 => (x"d8",x"87",x"eb",x"e5"),
  1221 => (x"66",x"c4",x"c1",x"86"),
  1222 => (x"01",x"a8",x"c0",x"48"),
  1223 => (x"a6",x"c8",x"87",x"c7"),
  1224 => (x"ce",x"78",x"c1",x"48"),
  1225 => (x"66",x"c4",x"c1",x"87"),
  1226 => (x"c8",x"88",x"c1",x"48"),
  1227 => (x"87",x"c3",x"58",x"a6"),
  1228 => (x"cc",x"87",x"f7",x"e4"),
  1229 => (x"78",x"c2",x"48",x"a6"),
  1230 => (x"cd",x"02",x"9c",x"74"),
  1231 => (x"66",x"c8",x"87",x"d6"),
  1232 => (x"66",x"c8",x"c1",x"48"),
  1233 => (x"cb",x"cd",x"03",x"a8"),
  1234 => (x"48",x"a6",x"d8",x"87"),
  1235 => (x"e9",x"e3",x"78",x"c0"),
  1236 => (x"c1",x"4c",x"70",x"87"),
  1237 => (x"c2",x"05",x"ac",x"d0"),
  1238 => (x"66",x"d8",x"87",x"d6"),
  1239 => (x"87",x"cd",x"e6",x"7e"),
  1240 => (x"a6",x"dc",x"49",x"70"),
  1241 => (x"87",x"d2",x"e3",x"59"),
  1242 => (x"ec",x"c0",x"4c",x"70"),
  1243 => (x"ea",x"c1",x"05",x"ac"),
  1244 => (x"49",x"66",x"c8",x"87"),
  1245 => (x"c0",x"c1",x"91",x"cb"),
  1246 => (x"a1",x"c4",x"81",x"66"),
  1247 => (x"c8",x"4d",x"6a",x"4a"),
  1248 => (x"66",x"d8",x"4a",x"a1"),
  1249 => (x"fc",x"c2",x"c1",x"52"),
  1250 => (x"87",x"ee",x"e2",x"79"),
  1251 => (x"02",x"9c",x"4c",x"70"),
  1252 => (x"fb",x"c0",x"87",x"d8"),
  1253 => (x"87",x"d2",x"02",x"ac"),
  1254 => (x"dd",x"e2",x"55",x"74"),
  1255 => (x"9c",x"4c",x"70",x"87"),
  1256 => (x"c0",x"87",x"c7",x"02"),
  1257 => (x"ff",x"05",x"ac",x"fb"),
  1258 => (x"e0",x"c0",x"87",x"ee"),
  1259 => (x"55",x"c1",x"c2",x"55"),
  1260 => (x"d4",x"7d",x"97",x"c0"),
  1261 => (x"a9",x"6e",x"49",x"66"),
  1262 => (x"c8",x"87",x"db",x"05"),
  1263 => (x"66",x"c4",x"48",x"66"),
  1264 => (x"87",x"ca",x"04",x"a8"),
  1265 => (x"c1",x"48",x"66",x"c8"),
  1266 => (x"58",x"a6",x"cc",x"80"),
  1267 => (x"66",x"c4",x"87",x"c8"),
  1268 => (x"c8",x"88",x"c1",x"48"),
  1269 => (x"e1",x"e1",x"58",x"a6"),
  1270 => (x"c1",x"4c",x"70",x"87"),
  1271 => (x"c8",x"05",x"ac",x"d0"),
  1272 => (x"48",x"66",x"d0",x"87"),
  1273 => (x"a6",x"d4",x"80",x"c1"),
  1274 => (x"ac",x"d0",x"c1",x"58"),
  1275 => (x"87",x"ea",x"fd",x"02"),
  1276 => (x"d4",x"48",x"a6",x"dc"),
  1277 => (x"66",x"d8",x"78",x"66"),
  1278 => (x"a8",x"66",x"dc",x"48"),
  1279 => (x"87",x"e6",x"c9",x"05"),
  1280 => (x"48",x"a6",x"e0",x"c0"),
  1281 => (x"c4",x"78",x"f0",x"c0"),
  1282 => (x"78",x"66",x"cc",x"80"),
  1283 => (x"78",x"c0",x"80",x"c4"),
  1284 => (x"c0",x"48",x"74",x"7e"),
  1285 => (x"f0",x"c0",x"88",x"fb"),
  1286 => (x"98",x"70",x"58",x"a6"),
  1287 => (x"87",x"e1",x"c8",x"02"),
  1288 => (x"c0",x"88",x"cb",x"48"),
  1289 => (x"70",x"58",x"a6",x"f0"),
  1290 => (x"e9",x"c0",x"02",x"98"),
  1291 => (x"88",x"c9",x"48",x"87"),
  1292 => (x"58",x"a6",x"f0",x"c0"),
  1293 => (x"c3",x"02",x"98",x"70"),
  1294 => (x"c4",x"48",x"87",x"e9"),
  1295 => (x"a6",x"f0",x"c0",x"88"),
  1296 => (x"02",x"98",x"70",x"58"),
  1297 => (x"c1",x"48",x"87",x"de"),
  1298 => (x"a6",x"f0",x"c0",x"88"),
  1299 => (x"02",x"98",x"70",x"58"),
  1300 => (x"c7",x"87",x"d0",x"c3"),
  1301 => (x"e0",x"c0",x"87",x"e5"),
  1302 => (x"78",x"c0",x"48",x"a6"),
  1303 => (x"c1",x"48",x"66",x"cc"),
  1304 => (x"58",x"a6",x"d0",x"80"),
  1305 => (x"87",x"d2",x"df",x"ff"),
  1306 => (x"ec",x"c0",x"4c",x"70"),
  1307 => (x"87",x"d7",x"02",x"ac"),
  1308 => (x"02",x"66",x"e0",x"c0"),
  1309 => (x"c0",x"87",x"c7",x"c0"),
  1310 => (x"c0",x"5c",x"a6",x"e4"),
  1311 => (x"48",x"74",x"87",x"c9"),
  1312 => (x"c0",x"88",x"f0",x"c0"),
  1313 => (x"c0",x"58",x"a6",x"e8"),
  1314 => (x"c0",x"02",x"ac",x"ec"),
  1315 => (x"de",x"ff",x"87",x"cd"),
  1316 => (x"4c",x"70",x"87",x"e8"),
  1317 => (x"05",x"ac",x"ec",x"c0"),
  1318 => (x"c0",x"87",x"f3",x"ff"),
  1319 => (x"d4",x"1e",x"66",x"e0"),
  1320 => (x"c0",x"1e",x"49",x"66"),
  1321 => (x"c1",x"1e",x"66",x"ec"),
  1322 => (x"d8",x"1e",x"e5",x"e2"),
  1323 => (x"fe",x"f4",x"49",x"66"),
  1324 => (x"ca",x"1e",x"c0",x"87"),
  1325 => (x"66",x"e0",x"c0",x"1e"),
  1326 => (x"c1",x"91",x"cb",x"49"),
  1327 => (x"d8",x"81",x"66",x"d8"),
  1328 => (x"a1",x"c4",x"48",x"a6"),
  1329 => (x"bf",x"66",x"d8",x"78"),
  1330 => (x"f1",x"de",x"ff",x"49"),
  1331 => (x"c0",x"86",x"d8",x"87"),
  1332 => (x"c1",x"06",x"a8",x"b7"),
  1333 => (x"1e",x"c1",x"87",x"c8"),
  1334 => (x"66",x"c8",x"1e",x"de"),
  1335 => (x"de",x"ff",x"49",x"bf"),
  1336 => (x"86",x"c8",x"87",x"dc"),
  1337 => (x"c0",x"48",x"49",x"70"),
  1338 => (x"e4",x"c0",x"88",x"08"),
  1339 => (x"b7",x"c0",x"58",x"a6"),
  1340 => (x"e9",x"c0",x"06",x"a8"),
  1341 => (x"66",x"e0",x"c0",x"87"),
  1342 => (x"a8",x"b7",x"dd",x"48"),
  1343 => (x"6e",x"87",x"df",x"03"),
  1344 => (x"e0",x"c0",x"49",x"bf"),
  1345 => (x"e0",x"c0",x"81",x"66"),
  1346 => (x"c1",x"49",x"66",x"51"),
  1347 => (x"81",x"bf",x"6e",x"81"),
  1348 => (x"c0",x"51",x"c1",x"c2"),
  1349 => (x"c2",x"49",x"66",x"e0"),
  1350 => (x"81",x"bf",x"6e",x"81"),
  1351 => (x"7e",x"c1",x"51",x"c0"),
  1352 => (x"ff",x"87",x"de",x"c4"),
  1353 => (x"c0",x"87",x"c6",x"df"),
  1354 => (x"ff",x"58",x"a6",x"e4"),
  1355 => (x"c0",x"87",x"fe",x"de"),
  1356 => (x"c0",x"58",x"a6",x"e8"),
  1357 => (x"c0",x"05",x"a8",x"ec"),
  1358 => (x"e4",x"c0",x"87",x"cb"),
  1359 => (x"e0",x"c0",x"48",x"a6"),
  1360 => (x"c4",x"c0",x"78",x"66"),
  1361 => (x"f1",x"db",x"ff",x"87"),
  1362 => (x"49",x"66",x"c8",x"87"),
  1363 => (x"c0",x"c1",x"91",x"cb"),
  1364 => (x"80",x"71",x"48",x"66"),
  1365 => (x"4a",x"6e",x"7e",x"70"),
  1366 => (x"49",x"6e",x"82",x"c8"),
  1367 => (x"e0",x"c0",x"81",x"ca"),
  1368 => (x"e4",x"c0",x"51",x"66"),
  1369 => (x"81",x"c1",x"49",x"66"),
  1370 => (x"89",x"66",x"e0",x"c0"),
  1371 => (x"30",x"71",x"48",x"c1"),
  1372 => (x"89",x"c1",x"49",x"70"),
  1373 => (x"c2",x"7a",x"97",x"71"),
  1374 => (x"49",x"bf",x"f5",x"ea"),
  1375 => (x"29",x"66",x"e0",x"c0"),
  1376 => (x"48",x"4a",x"6a",x"97"),
  1377 => (x"f0",x"c0",x"98",x"71"),
  1378 => (x"49",x"6e",x"58",x"a6"),
  1379 => (x"4d",x"69",x"81",x"c4"),
  1380 => (x"d8",x"48",x"66",x"dc"),
  1381 => (x"c0",x"02",x"a8",x"66"),
  1382 => (x"a6",x"d8",x"87",x"c8"),
  1383 => (x"c0",x"78",x"c0",x"48"),
  1384 => (x"a6",x"d8",x"87",x"c5"),
  1385 => (x"d8",x"78",x"c1",x"48"),
  1386 => (x"e0",x"c0",x"1e",x"66"),
  1387 => (x"ff",x"49",x"75",x"1e"),
  1388 => (x"c8",x"87",x"cb",x"db"),
  1389 => (x"c0",x"4c",x"70",x"86"),
  1390 => (x"c1",x"06",x"ac",x"b7"),
  1391 => (x"85",x"74",x"87",x"d4"),
  1392 => (x"74",x"49",x"e0",x"c0"),
  1393 => (x"c1",x"4b",x"75",x"89"),
  1394 => (x"71",x"4a",x"ed",x"db"),
  1395 => (x"87",x"d8",x"eb",x"fe"),
  1396 => (x"e8",x"c0",x"85",x"c2"),
  1397 => (x"80",x"c1",x"48",x"66"),
  1398 => (x"58",x"a6",x"ec",x"c0"),
  1399 => (x"49",x"66",x"ec",x"c0"),
  1400 => (x"a9",x"70",x"81",x"c1"),
  1401 => (x"87",x"c8",x"c0",x"02"),
  1402 => (x"c0",x"48",x"a6",x"d8"),
  1403 => (x"87",x"c5",x"c0",x"78"),
  1404 => (x"c1",x"48",x"a6",x"d8"),
  1405 => (x"1e",x"66",x"d8",x"78"),
  1406 => (x"c0",x"49",x"a4",x"c2"),
  1407 => (x"88",x"71",x"48",x"e0"),
  1408 => (x"75",x"1e",x"49",x"70"),
  1409 => (x"f5",x"d9",x"ff",x"49"),
  1410 => (x"c0",x"86",x"c8",x"87"),
  1411 => (x"ff",x"01",x"a8",x"b7"),
  1412 => (x"e8",x"c0",x"87",x"c0"),
  1413 => (x"d1",x"c0",x"02",x"66"),
  1414 => (x"c9",x"49",x"6e",x"87"),
  1415 => (x"66",x"e8",x"c0",x"81"),
  1416 => (x"c1",x"48",x"6e",x"51"),
  1417 => (x"c0",x"78",x"cc",x"c4"),
  1418 => (x"49",x"6e",x"87",x"cc"),
  1419 => (x"51",x"c2",x"81",x"c9"),
  1420 => (x"c5",x"c1",x"48",x"6e"),
  1421 => (x"7e",x"c1",x"78",x"c0"),
  1422 => (x"ff",x"87",x"c6",x"c0"),
  1423 => (x"70",x"87",x"eb",x"d8"),
  1424 => (x"c0",x"02",x"6e",x"4c"),
  1425 => (x"66",x"c8",x"87",x"f5"),
  1426 => (x"a8",x"66",x"c4",x"48"),
  1427 => (x"87",x"cb",x"c0",x"04"),
  1428 => (x"c1",x"48",x"66",x"c8"),
  1429 => (x"58",x"a6",x"cc",x"80"),
  1430 => (x"c4",x"87",x"e0",x"c0"),
  1431 => (x"88",x"c1",x"48",x"66"),
  1432 => (x"c0",x"58",x"a6",x"c8"),
  1433 => (x"c6",x"c1",x"87",x"d5"),
  1434 => (x"c8",x"c0",x"05",x"ac"),
  1435 => (x"48",x"66",x"cc",x"87"),
  1436 => (x"a6",x"d0",x"80",x"c1"),
  1437 => (x"f1",x"d7",x"ff",x"58"),
  1438 => (x"d0",x"4c",x"70",x"87"),
  1439 => (x"80",x"c1",x"48",x"66"),
  1440 => (x"74",x"58",x"a6",x"d4"),
  1441 => (x"cb",x"c0",x"02",x"9c"),
  1442 => (x"48",x"66",x"c8",x"87"),
  1443 => (x"a8",x"66",x"c8",x"c1"),
  1444 => (x"87",x"f5",x"f2",x"04"),
  1445 => (x"87",x"c9",x"d7",x"ff"),
  1446 => (x"c7",x"48",x"66",x"c8"),
  1447 => (x"e5",x"c0",x"03",x"a8"),
  1448 => (x"c8",x"e7",x"c2",x"87"),
  1449 => (x"c8",x"78",x"c0",x"48"),
  1450 => (x"91",x"cb",x"49",x"66"),
  1451 => (x"81",x"66",x"c0",x"c1"),
  1452 => (x"6a",x"4a",x"a1",x"c4"),
  1453 => (x"79",x"52",x"c0",x"4a"),
  1454 => (x"c1",x"48",x"66",x"c8"),
  1455 => (x"58",x"a6",x"cc",x"80"),
  1456 => (x"ff",x"04",x"a8",x"c7"),
  1457 => (x"d0",x"ff",x"87",x"db"),
  1458 => (x"e9",x"de",x"ff",x"8e"),
  1459 => (x"61",x"6f",x"4c",x"87"),
  1460 => (x"65",x"53",x"20",x"64"),
  1461 => (x"6e",x"69",x"74",x"74"),
  1462 => (x"81",x"20",x"73",x"67"),
  1463 => (x"76",x"61",x"53",x"00"),
  1464 => (x"65",x"53",x"20",x"65"),
  1465 => (x"6e",x"69",x"74",x"74"),
  1466 => (x"81",x"20",x"73",x"67"),
  1467 => (x"00",x"20",x"3a",x"00"),
  1468 => (x"71",x"1e",x"73",x"1e"),
  1469 => (x"c6",x"02",x"9b",x"4b"),
  1470 => (x"c4",x"e7",x"c2",x"87"),
  1471 => (x"c7",x"78",x"c0",x"48"),
  1472 => (x"c4",x"e7",x"c2",x"1e"),
  1473 => (x"c1",x"1e",x"49",x"bf"),
  1474 => (x"c2",x"1e",x"f2",x"e0"),
  1475 => (x"49",x"bf",x"c0",x"e7"),
  1476 => (x"cc",x"87",x"d1",x"ec"),
  1477 => (x"c0",x"e7",x"c2",x"86"),
  1478 => (x"c7",x"e7",x"49",x"bf"),
  1479 => (x"02",x"9b",x"73",x"87"),
  1480 => (x"e0",x"c1",x"87",x"c8"),
  1481 => (x"e6",x"c0",x"49",x"f2"),
  1482 => (x"dd",x"ff",x"87",x"e5"),
  1483 => (x"73",x"1e",x"87",x"cc"),
  1484 => (x"c1",x"4b",x"c0",x"1e"),
  1485 => (x"c0",x"49",x"d9",x"dd"),
  1486 => (x"c2",x"87",x"ff",x"fa"),
  1487 => (x"c0",x"48",x"fa",x"d5"),
  1488 => (x"d5",x"e2",x"c1",x"50"),
  1489 => (x"f4",x"c0",x"49",x"bf"),
  1490 => (x"98",x"70",x"87",x"d5"),
  1491 => (x"c1",x"87",x"c4",x"05"),
  1492 => (x"73",x"4b",x"e5",x"dd"),
  1493 => (x"e1",x"dc",x"ff",x"48"),
  1494 => (x"43",x"49",x"56",x"87"),
  1495 => (x"20",x"20",x"30",x"32"),
  1496 => (x"47",x"46",x"43",x"20"),
  1497 => (x"4d",x"4f",x"52",x"00"),
  1498 => (x"61",x"6f",x"6c",x"20"),
  1499 => (x"67",x"6e",x"69",x"64"),
  1500 => (x"69",x"61",x"66",x"20"),
  1501 => (x"00",x"64",x"65",x"6c"),
  1502 => (x"87",x"c8",x"c8",x"1e"),
  1503 => (x"ef",x"fd",x"49",x"c1"),
  1504 => (x"f6",x"ec",x"fe",x"87"),
  1505 => (x"02",x"98",x"70",x"87"),
  1506 => (x"f5",x"fe",x"87",x"cd"),
  1507 => (x"98",x"70",x"87",x"f3"),
  1508 => (x"c1",x"87",x"c4",x"02"),
  1509 => (x"c0",x"87",x"c2",x"4a"),
  1510 => (x"05",x"9a",x"72",x"4a"),
  1511 => (x"1e",x"c0",x"87",x"ce"),
  1512 => (x"49",x"cc",x"df",x"c1"),
  1513 => (x"87",x"f5",x"f0",x"c0"),
  1514 => (x"87",x"fe",x"86",x"c4"),
  1515 => (x"87",x"f4",x"f7",x"c0"),
  1516 => (x"df",x"c1",x"1e",x"c0"),
  1517 => (x"f0",x"c0",x"49",x"d7"),
  1518 => (x"1e",x"c0",x"87",x"e3"),
  1519 => (x"70",x"87",x"ef",x"fd"),
  1520 => (x"d8",x"f0",x"c0",x"49"),
  1521 => (x"87",x"fb",x"c3",x"87"),
  1522 => (x"4f",x"26",x"8e",x"f8"),
  1523 => (x"66",x"20",x"44",x"53"),
  1524 => (x"65",x"6c",x"69",x"61"),
  1525 => (x"42",x"00",x"2e",x"64"),
  1526 => (x"69",x"74",x"6f",x"6f"),
  1527 => (x"2e",x"2e",x"67",x"6e"),
  1528 => (x"c0",x"1e",x"00",x"2e"),
  1529 => (x"fa",x"87",x"c4",x"e8"),
  1530 => (x"1e",x"4f",x"26",x"87"),
  1531 => (x"48",x"c4",x"e7",x"c2"),
  1532 => (x"e7",x"c2",x"78",x"c0"),
  1533 => (x"78",x"c0",x"48",x"c0"),
  1534 => (x"e5",x"87",x"fd",x"fd"),
  1535 => (x"26",x"48",x"c0",x"87"),
  1536 => (x"20",x"20",x"20",x"4f"),
  1537 => (x"20",x"20",x"20",x"20"),
  1538 => (x"20",x"20",x"20",x"20"),
  1539 => (x"78",x"45",x"20",x"20"),
  1540 => (x"20",x"20",x"74",x"69"),
  1541 => (x"20",x"20",x"20",x"20"),
  1542 => (x"20",x"20",x"20",x"20"),
  1543 => (x"00",x"81",x"20",x"20"),
  1544 => (x"20",x"20",x"20",x"80"),
  1545 => (x"20",x"20",x"20",x"20"),
  1546 => (x"20",x"20",x"20",x"20"),
  1547 => (x"63",x"61",x"42",x"20"),
  1548 => (x"10",x"bc",x"00",x"6b"),
  1549 => (x"29",x"d9",x"00",x"00"),
  1550 => (x"00",x"00",x"00",x"00"),
  1551 => (x"00",x"10",x"bc",x"00"),
  1552 => (x"00",x"29",x"f7",x"00"),
  1553 => (x"00",x"00",x"00",x"00"),
  1554 => (x"00",x"00",x"10",x"bc"),
  1555 => (x"00",x"00",x"2a",x"15"),
  1556 => (x"bc",x"00",x"00",x"00"),
  1557 => (x"33",x"00",x"00",x"10"),
  1558 => (x"00",x"00",x"00",x"2a"),
  1559 => (x"10",x"bc",x"00",x"00"),
  1560 => (x"2a",x"51",x"00",x"00"),
  1561 => (x"00",x"00",x"00",x"00"),
  1562 => (x"00",x"10",x"bc",x"00"),
  1563 => (x"00",x"2a",x"6f",x"00"),
  1564 => (x"00",x"00",x"00",x"00"),
  1565 => (x"00",x"00",x"10",x"bc"),
  1566 => (x"00",x"00",x"2a",x"8d"),
  1567 => (x"bc",x"00",x"00",x"00"),
  1568 => (x"00",x"00",x"00",x"10"),
  1569 => (x"00",x"00",x"00",x"00"),
  1570 => (x"11",x"51",x"00",x"00"),
  1571 => (x"00",x"00",x"00",x"00"),
  1572 => (x"00",x"00",x"00",x"00"),
  1573 => (x"00",x"18",x"99",x"00"),
  1574 => (x"43",x"49",x"56",x"00"),
  1575 => (x"20",x"20",x"30",x"32"),
  1576 => (x"4d",x"4f",x"52",x"20"),
  1577 => (x"61",x"6f",x"4c",x"00"),
  1578 => (x"2e",x"2a",x"20",x"64"),
  1579 => (x"f0",x"fe",x"1e",x"00"),
  1580 => (x"cd",x"78",x"c0",x"48"),
  1581 => (x"26",x"09",x"79",x"09"),
  1582 => (x"fe",x"1e",x"1e",x"4f"),
  1583 => (x"48",x"7e",x"bf",x"f0"),
  1584 => (x"1e",x"4f",x"26",x"26"),
  1585 => (x"c1",x"48",x"f0",x"fe"),
  1586 => (x"1e",x"4f",x"26",x"78"),
  1587 => (x"c0",x"48",x"f0",x"fe"),
  1588 => (x"1e",x"4f",x"26",x"78"),
  1589 => (x"52",x"c0",x"4a",x"71"),
  1590 => (x"0e",x"4f",x"26",x"52"),
  1591 => (x"5d",x"5c",x"5b",x"5e"),
  1592 => (x"71",x"86",x"f4",x"0e"),
  1593 => (x"7e",x"6d",x"97",x"4d"),
  1594 => (x"97",x"4c",x"a5",x"c1"),
  1595 => (x"a6",x"c8",x"48",x"6c"),
  1596 => (x"c4",x"48",x"6e",x"58"),
  1597 => (x"c5",x"05",x"a8",x"66"),
  1598 => (x"c0",x"48",x"ff",x"87"),
  1599 => (x"ca",x"ff",x"87",x"e6"),
  1600 => (x"49",x"a5",x"c2",x"87"),
  1601 => (x"71",x"4b",x"6c",x"97"),
  1602 => (x"6b",x"97",x"4b",x"a3"),
  1603 => (x"7e",x"6c",x"97",x"4b"),
  1604 => (x"80",x"c1",x"48",x"6e"),
  1605 => (x"c7",x"58",x"a6",x"c8"),
  1606 => (x"58",x"a6",x"cc",x"98"),
  1607 => (x"fe",x"7c",x"97",x"70"),
  1608 => (x"48",x"73",x"87",x"e1"),
  1609 => (x"4d",x"26",x"8e",x"f4"),
  1610 => (x"4b",x"26",x"4c",x"26"),
  1611 => (x"5e",x"0e",x"4f",x"26"),
  1612 => (x"f4",x"0e",x"5c",x"5b"),
  1613 => (x"d8",x"4c",x"71",x"86"),
  1614 => (x"ff",x"c3",x"4a",x"66"),
  1615 => (x"4b",x"a4",x"c2",x"9a"),
  1616 => (x"73",x"49",x"6c",x"97"),
  1617 => (x"51",x"72",x"49",x"a1"),
  1618 => (x"6e",x"7e",x"6c",x"97"),
  1619 => (x"c8",x"80",x"c1",x"48"),
  1620 => (x"98",x"c7",x"58",x"a6"),
  1621 => (x"70",x"58",x"a6",x"cc"),
  1622 => (x"ff",x"8e",x"f4",x"54"),
  1623 => (x"1e",x"1e",x"87",x"ca"),
  1624 => (x"e0",x"87",x"e8",x"fd"),
  1625 => (x"c0",x"49",x"4a",x"bf"),
  1626 => (x"02",x"99",x"c0",x"e0"),
  1627 => (x"1e",x"72",x"87",x"cb"),
  1628 => (x"49",x"eb",x"ea",x"c2"),
  1629 => (x"c4",x"87",x"f7",x"fe"),
  1630 => (x"87",x"fd",x"fc",x"86"),
  1631 => (x"c2",x"fd",x"7e",x"70"),
  1632 => (x"4f",x"26",x"26",x"87"),
  1633 => (x"eb",x"ea",x"c2",x"1e"),
  1634 => (x"87",x"c7",x"fd",x"49"),
  1635 => (x"49",x"de",x"e5",x"c1"),
  1636 => (x"c5",x"87",x"da",x"fc"),
  1637 => (x"4f",x"26",x"87",x"d9"),
  1638 => (x"5c",x"5b",x"5e",x"0e"),
  1639 => (x"eb",x"c2",x"0e",x"5d"),
  1640 => (x"c1",x"4a",x"bf",x"ca"),
  1641 => (x"49",x"bf",x"ec",x"e7"),
  1642 => (x"71",x"bc",x"72",x"4c"),
  1643 => (x"87",x"db",x"fc",x"4d"),
  1644 => (x"49",x"74",x"4b",x"c0"),
  1645 => (x"d5",x"02",x"99",x"d0"),
  1646 => (x"d0",x"49",x"75",x"87"),
  1647 => (x"c0",x"1e",x"71",x"99"),
  1648 => (x"fe",x"ed",x"c1",x"1e"),
  1649 => (x"12",x"82",x"73",x"4a"),
  1650 => (x"87",x"e4",x"c0",x"49"),
  1651 => (x"2c",x"c1",x"86",x"c8"),
  1652 => (x"ab",x"c8",x"83",x"2d"),
  1653 => (x"87",x"da",x"ff",x"04"),
  1654 => (x"c1",x"87",x"e8",x"fb"),
  1655 => (x"c2",x"48",x"ec",x"e7"),
  1656 => (x"78",x"bf",x"ca",x"eb"),
  1657 => (x"4c",x"26",x"4d",x"26"),
  1658 => (x"4f",x"26",x"4b",x"26"),
  1659 => (x"00",x"00",x"00",x"00"),
  1660 => (x"48",x"d0",x"ff",x"1e"),
  1661 => (x"ff",x"78",x"e1",x"c8"),
  1662 => (x"78",x"c5",x"48",x"d4"),
  1663 => (x"c3",x"02",x"66",x"c4"),
  1664 => (x"78",x"e0",x"c3",x"87"),
  1665 => (x"c6",x"02",x"66",x"c8"),
  1666 => (x"48",x"d4",x"ff",x"87"),
  1667 => (x"ff",x"78",x"f0",x"c3"),
  1668 => (x"78",x"71",x"48",x"d4"),
  1669 => (x"c8",x"48",x"d0",x"ff"),
  1670 => (x"e0",x"c0",x"78",x"e1"),
  1671 => (x"0e",x"4f",x"26",x"78"),
  1672 => (x"0e",x"5c",x"5b",x"5e"),
  1673 => (x"ea",x"c2",x"4c",x"71"),
  1674 => (x"ee",x"fa",x"49",x"eb"),
  1675 => (x"c0",x"4a",x"70",x"87"),
  1676 => (x"c2",x"04",x"aa",x"b7"),
  1677 => (x"e0",x"c3",x"87",x"e3"),
  1678 => (x"87",x"c9",x"05",x"aa"),
  1679 => (x"48",x"e2",x"eb",x"c1"),
  1680 => (x"d4",x"c2",x"78",x"c1"),
  1681 => (x"aa",x"f0",x"c3",x"87"),
  1682 => (x"c1",x"87",x"c9",x"05"),
  1683 => (x"c1",x"48",x"de",x"eb"),
  1684 => (x"87",x"f5",x"c1",x"78"),
  1685 => (x"bf",x"e2",x"eb",x"c1"),
  1686 => (x"72",x"87",x"c7",x"02"),
  1687 => (x"b3",x"c0",x"c2",x"4b"),
  1688 => (x"4b",x"72",x"87",x"c2"),
  1689 => (x"d1",x"05",x"9c",x"74"),
  1690 => (x"de",x"eb",x"c1",x"87"),
  1691 => (x"eb",x"c1",x"1e",x"bf"),
  1692 => (x"72",x"1e",x"bf",x"e2"),
  1693 => (x"87",x"f8",x"fd",x"49"),
  1694 => (x"eb",x"c1",x"86",x"c8"),
  1695 => (x"c0",x"02",x"bf",x"de"),
  1696 => (x"49",x"73",x"87",x"e0"),
  1697 => (x"91",x"29",x"b7",x"c4"),
  1698 => (x"81",x"fe",x"ec",x"c1"),
  1699 => (x"9a",x"cf",x"4a",x"73"),
  1700 => (x"48",x"c1",x"92",x"c2"),
  1701 => (x"4a",x"70",x"30",x"72"),
  1702 => (x"48",x"72",x"ba",x"ff"),
  1703 => (x"79",x"70",x"98",x"69"),
  1704 => (x"49",x"73",x"87",x"db"),
  1705 => (x"91",x"29",x"b7",x"c4"),
  1706 => (x"81",x"fe",x"ec",x"c1"),
  1707 => (x"9a",x"cf",x"4a",x"73"),
  1708 => (x"48",x"c3",x"92",x"c2"),
  1709 => (x"4a",x"70",x"30",x"72"),
  1710 => (x"70",x"b0",x"69",x"48"),
  1711 => (x"e2",x"eb",x"c1",x"79"),
  1712 => (x"c1",x"78",x"c0",x"48"),
  1713 => (x"c0",x"48",x"de",x"eb"),
  1714 => (x"eb",x"ea",x"c2",x"78"),
  1715 => (x"87",x"cb",x"f8",x"49"),
  1716 => (x"b7",x"c0",x"4a",x"70"),
  1717 => (x"dd",x"fd",x"03",x"aa"),
  1718 => (x"fc",x"48",x"c0",x"87"),
  1719 => (x"00",x"00",x"87",x"c8"),
  1720 => (x"00",x"00",x"00",x"00"),
  1721 => (x"71",x"1e",x"00",x"00"),
  1722 => (x"f2",x"fc",x"49",x"4a"),
  1723 => (x"1e",x"4f",x"26",x"87"),
  1724 => (x"49",x"72",x"4a",x"c0"),
  1725 => (x"ec",x"c1",x"91",x"c4"),
  1726 => (x"79",x"c0",x"81",x"fe"),
  1727 => (x"b7",x"d0",x"82",x"c1"),
  1728 => (x"87",x"ee",x"04",x"aa"),
  1729 => (x"5e",x"0e",x"4f",x"26"),
  1730 => (x"0e",x"5d",x"5c",x"5b"),
  1731 => (x"fa",x"f6",x"4d",x"71"),
  1732 => (x"c4",x"4a",x"75",x"87"),
  1733 => (x"c1",x"92",x"2a",x"b7"),
  1734 => (x"75",x"82",x"fe",x"ec"),
  1735 => (x"c2",x"9c",x"cf",x"4c"),
  1736 => (x"4b",x"49",x"6a",x"94"),
  1737 => (x"9b",x"c3",x"2b",x"74"),
  1738 => (x"30",x"74",x"48",x"c2"),
  1739 => (x"bc",x"ff",x"4c",x"70"),
  1740 => (x"98",x"71",x"48",x"74"),
  1741 => (x"ca",x"f6",x"7a",x"70"),
  1742 => (x"fa",x"48",x"73",x"87"),
  1743 => (x"00",x"00",x"87",x"e6"),
  1744 => (x"00",x"00",x"00",x"00"),
  1745 => (x"00",x"00",x"00",x"00"),
  1746 => (x"00",x"00",x"00",x"00"),
  1747 => (x"00",x"00",x"00",x"00"),
  1748 => (x"00",x"00",x"00",x"00"),
  1749 => (x"00",x"00",x"00",x"00"),
  1750 => (x"00",x"00",x"00",x"00"),
  1751 => (x"00",x"00",x"00",x"00"),
  1752 => (x"00",x"00",x"00",x"00"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"00",x"00",x"00"),
  1755 => (x"00",x"00",x"00",x"00"),
  1756 => (x"00",x"00",x"00",x"00"),
  1757 => (x"00",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"00",x"00"),
  1759 => (x"1e",x"16",x"00",x"00"),
  1760 => (x"36",x"2e",x"25",x"26"),
  1761 => (x"ff",x"1e",x"3e",x"3d"),
  1762 => (x"e1",x"c8",x"48",x"d0"),
  1763 => (x"ff",x"48",x"71",x"78"),
  1764 => (x"c4",x"78",x"08",x"d4"),
  1765 => (x"d4",x"ff",x"48",x"66"),
  1766 => (x"4f",x"26",x"78",x"08"),
  1767 => (x"c4",x"4a",x"71",x"1e"),
  1768 => (x"e0",x"c1",x"1e",x"66"),
  1769 => (x"dd",x"ff",x"49",x"a2"),
  1770 => (x"49",x"66",x"c8",x"87"),
  1771 => (x"ff",x"29",x"b7",x"c8"),
  1772 => (x"78",x"71",x"48",x"d4"),
  1773 => (x"c0",x"48",x"d0",x"ff"),
  1774 => (x"26",x"26",x"78",x"e0"),
  1775 => (x"d4",x"ff",x"1e",x"4f"),
  1776 => (x"7a",x"ff",x"c3",x"4a"),
  1777 => (x"c8",x"48",x"d0",x"ff"),
  1778 => (x"7a",x"de",x"78",x"e1"),
  1779 => (x"bf",x"f5",x"ea",x"c2"),
  1780 => (x"c8",x"48",x"49",x"7a"),
  1781 => (x"71",x"7a",x"70",x"28"),
  1782 => (x"70",x"28",x"d0",x"48"),
  1783 => (x"d8",x"48",x"71",x"7a"),
  1784 => (x"ff",x"7a",x"70",x"28"),
  1785 => (x"e0",x"c0",x"48",x"d0"),
  1786 => (x"0e",x"4f",x"26",x"78"),
  1787 => (x"5d",x"5c",x"5b",x"5e"),
  1788 => (x"c2",x"4c",x"71",x"0e"),
  1789 => (x"4d",x"bf",x"f5",x"ea"),
  1790 => (x"d0",x"2b",x"74",x"4b"),
  1791 => (x"83",x"c1",x"9b",x"66"),
  1792 => (x"04",x"ab",x"66",x"d4"),
  1793 => (x"4b",x"c0",x"87",x"c2"),
  1794 => (x"66",x"d0",x"4a",x"74"),
  1795 => (x"ff",x"31",x"72",x"49"),
  1796 => (x"73",x"99",x"75",x"b9"),
  1797 => (x"70",x"30",x"72",x"48"),
  1798 => (x"b0",x"71",x"48",x"4a"),
  1799 => (x"58",x"f9",x"ea",x"c2"),
  1800 => (x"26",x"87",x"da",x"fe"),
  1801 => (x"26",x"4c",x"26",x"4d"),
  1802 => (x"1e",x"4f",x"26",x"4b"),
  1803 => (x"c8",x"48",x"d0",x"ff"),
  1804 => (x"48",x"71",x"78",x"c9"),
  1805 => (x"78",x"08",x"d4",x"ff"),
  1806 => (x"71",x"1e",x"4f",x"26"),
  1807 => (x"87",x"eb",x"49",x"4a"),
  1808 => (x"c8",x"48",x"d0",x"ff"),
  1809 => (x"1e",x"4f",x"26",x"78"),
  1810 => (x"4b",x"71",x"1e",x"73"),
  1811 => (x"bf",x"c5",x"eb",x"c2"),
  1812 => (x"c2",x"87",x"c3",x"02"),
  1813 => (x"d0",x"ff",x"87",x"eb"),
  1814 => (x"78",x"c9",x"c8",x"48"),
  1815 => (x"e0",x"c0",x"49",x"73"),
  1816 => (x"48",x"d4",x"ff",x"b1"),
  1817 => (x"ea",x"c2",x"78",x"71"),
  1818 => (x"78",x"c0",x"48",x"f9"),
  1819 => (x"c5",x"02",x"66",x"c8"),
  1820 => (x"49",x"ff",x"c3",x"87"),
  1821 => (x"49",x"c0",x"87",x"c2"),
  1822 => (x"59",x"c1",x"eb",x"c2"),
  1823 => (x"c6",x"02",x"66",x"cc"),
  1824 => (x"d5",x"d5",x"c5",x"87"),
  1825 => (x"cf",x"87",x"c4",x"4a"),
  1826 => (x"c2",x"4a",x"ff",x"ff"),
  1827 => (x"c2",x"5a",x"c5",x"eb"),
  1828 => (x"c1",x"48",x"c5",x"eb"),
  1829 => (x"26",x"87",x"c4",x"78"),
  1830 => (x"26",x"4c",x"26",x"4d"),
  1831 => (x"0e",x"4f",x"26",x"4b"),
  1832 => (x"5d",x"5c",x"5b",x"5e"),
  1833 => (x"c2",x"4a",x"71",x"0e"),
  1834 => (x"4c",x"bf",x"c1",x"eb"),
  1835 => (x"cb",x"02",x"9a",x"72"),
  1836 => (x"91",x"c8",x"49",x"87"),
  1837 => (x"4b",x"fd",x"f0",x"c1"),
  1838 => (x"87",x"c4",x"83",x"71"),
  1839 => (x"4b",x"fd",x"f4",x"c1"),
  1840 => (x"49",x"13",x"4d",x"c0"),
  1841 => (x"ea",x"c2",x"99",x"74"),
  1842 => (x"ff",x"b9",x"bf",x"fd"),
  1843 => (x"78",x"71",x"48",x"d4"),
  1844 => (x"85",x"2c",x"b7",x"c1"),
  1845 => (x"04",x"ad",x"b7",x"c8"),
  1846 => (x"ea",x"c2",x"87",x"e8"),
  1847 => (x"c8",x"48",x"bf",x"f9"),
  1848 => (x"fd",x"ea",x"c2",x"80"),
  1849 => (x"87",x"ef",x"fe",x"58"),
  1850 => (x"71",x"1e",x"73",x"1e"),
  1851 => (x"9a",x"4a",x"13",x"4b"),
  1852 => (x"72",x"87",x"cb",x"02"),
  1853 => (x"87",x"e7",x"fe",x"49"),
  1854 => (x"05",x"9a",x"4a",x"13"),
  1855 => (x"da",x"fe",x"87",x"f5"),
  1856 => (x"ea",x"c2",x"1e",x"87"),
  1857 => (x"c2",x"49",x"bf",x"f9"),
  1858 => (x"c1",x"48",x"f9",x"ea"),
  1859 => (x"c0",x"c4",x"78",x"a1"),
  1860 => (x"db",x"03",x"a9",x"b7"),
  1861 => (x"48",x"d4",x"ff",x"87"),
  1862 => (x"bf",x"fd",x"ea",x"c2"),
  1863 => (x"f9",x"ea",x"c2",x"78"),
  1864 => (x"ea",x"c2",x"49",x"bf"),
  1865 => (x"a1",x"c1",x"48",x"f9"),
  1866 => (x"b7",x"c0",x"c4",x"78"),
  1867 => (x"87",x"e5",x"04",x"a9"),
  1868 => (x"c8",x"48",x"d0",x"ff"),
  1869 => (x"c5",x"eb",x"c2",x"78"),
  1870 => (x"26",x"78",x"c0",x"48"),
  1871 => (x"00",x"00",x"00",x"4f"),
  1872 => (x"00",x"00",x"00",x"00"),
  1873 => (x"00",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"5f",x"5f"),
  1875 => (x"03",x"03",x"00",x"00"),
  1876 => (x"00",x"03",x"03",x"00"),
  1877 => (x"7f",x"7f",x"14",x"00"),
  1878 => (x"14",x"7f",x"7f",x"14"),
  1879 => (x"2e",x"24",x"00",x"00"),
  1880 => (x"12",x"3a",x"6b",x"6b"),
  1881 => (x"36",x"6a",x"4c",x"00"),
  1882 => (x"32",x"56",x"6c",x"18"),
  1883 => (x"4f",x"7e",x"30",x"00"),
  1884 => (x"68",x"3a",x"77",x"59"),
  1885 => (x"04",x"00",x"00",x"40"),
  1886 => (x"00",x"00",x"03",x"07"),
  1887 => (x"1c",x"00",x"00",x"00"),
  1888 => (x"00",x"41",x"63",x"3e"),
  1889 => (x"41",x"00",x"00",x"00"),
  1890 => (x"00",x"1c",x"3e",x"63"),
  1891 => (x"3e",x"2a",x"08",x"00"),
  1892 => (x"2a",x"3e",x"1c",x"1c"),
  1893 => (x"08",x"08",x"00",x"08"),
  1894 => (x"08",x"08",x"3e",x"3e"),
  1895 => (x"80",x"00",x"00",x"00"),
  1896 => (x"00",x"00",x"60",x"e0"),
  1897 => (x"08",x"08",x"00",x"00"),
  1898 => (x"08",x"08",x"08",x"08"),
  1899 => (x"00",x"00",x"00",x"00"),
  1900 => (x"00",x"00",x"60",x"60"),
  1901 => (x"30",x"60",x"40",x"00"),
  1902 => (x"03",x"06",x"0c",x"18"),
  1903 => (x"7f",x"3e",x"00",x"01"),
  1904 => (x"3e",x"7f",x"4d",x"59"),
  1905 => (x"06",x"04",x"00",x"00"),
  1906 => (x"00",x"00",x"7f",x"7f"),
  1907 => (x"63",x"42",x"00",x"00"),
  1908 => (x"46",x"4f",x"59",x"71"),
  1909 => (x"63",x"22",x"00",x"00"),
  1910 => (x"36",x"7f",x"49",x"49"),
  1911 => (x"16",x"1c",x"18",x"00"),
  1912 => (x"10",x"7f",x"7f",x"13"),
  1913 => (x"67",x"27",x"00",x"00"),
  1914 => (x"39",x"7d",x"45",x"45"),
  1915 => (x"7e",x"3c",x"00",x"00"),
  1916 => (x"30",x"79",x"49",x"4b"),
  1917 => (x"01",x"01",x"00",x"00"),
  1918 => (x"07",x"0f",x"79",x"71"),
  1919 => (x"7f",x"36",x"00",x"00"),
  1920 => (x"36",x"7f",x"49",x"49"),
  1921 => (x"4f",x"06",x"00",x"00"),
  1922 => (x"1e",x"3f",x"69",x"49"),
  1923 => (x"00",x"00",x"00",x"00"),
  1924 => (x"00",x"00",x"66",x"66"),
  1925 => (x"80",x"00",x"00",x"00"),
  1926 => (x"00",x"00",x"66",x"e6"),
  1927 => (x"08",x"08",x"00",x"00"),
  1928 => (x"22",x"22",x"14",x"14"),
  1929 => (x"14",x"14",x"00",x"00"),
  1930 => (x"14",x"14",x"14",x"14"),
  1931 => (x"22",x"22",x"00",x"00"),
  1932 => (x"08",x"08",x"14",x"14"),
  1933 => (x"03",x"02",x"00",x"00"),
  1934 => (x"06",x"0f",x"59",x"51"),
  1935 => (x"41",x"7f",x"3e",x"00"),
  1936 => (x"1e",x"1f",x"55",x"5d"),
  1937 => (x"7f",x"7e",x"00",x"00"),
  1938 => (x"7e",x"7f",x"09",x"09"),
  1939 => (x"7f",x"7f",x"00",x"00"),
  1940 => (x"36",x"7f",x"49",x"49"),
  1941 => (x"3e",x"1c",x"00",x"00"),
  1942 => (x"41",x"41",x"41",x"63"),
  1943 => (x"7f",x"7f",x"00",x"00"),
  1944 => (x"1c",x"3e",x"63",x"41"),
  1945 => (x"7f",x"7f",x"00",x"00"),
  1946 => (x"41",x"41",x"49",x"49"),
  1947 => (x"7f",x"7f",x"00",x"00"),
  1948 => (x"01",x"01",x"09",x"09"),
  1949 => (x"7f",x"3e",x"00",x"00"),
  1950 => (x"7a",x"7b",x"49",x"41"),
  1951 => (x"7f",x"7f",x"00",x"00"),
  1952 => (x"7f",x"7f",x"08",x"08"),
  1953 => (x"41",x"00",x"00",x"00"),
  1954 => (x"00",x"41",x"7f",x"7f"),
  1955 => (x"60",x"20",x"00",x"00"),
  1956 => (x"3f",x"7f",x"40",x"40"),
  1957 => (x"08",x"7f",x"7f",x"00"),
  1958 => (x"41",x"63",x"36",x"1c"),
  1959 => (x"7f",x"7f",x"00",x"00"),
  1960 => (x"40",x"40",x"40",x"40"),
  1961 => (x"06",x"7f",x"7f",x"00"),
  1962 => (x"7f",x"7f",x"06",x"0c"),
  1963 => (x"06",x"7f",x"7f",x"00"),
  1964 => (x"7f",x"7f",x"18",x"0c"),
  1965 => (x"7f",x"3e",x"00",x"00"),
  1966 => (x"3e",x"7f",x"41",x"41"),
  1967 => (x"7f",x"7f",x"00",x"00"),
  1968 => (x"06",x"0f",x"09",x"09"),
  1969 => (x"41",x"7f",x"3e",x"00"),
  1970 => (x"40",x"7e",x"7f",x"61"),
  1971 => (x"7f",x"7f",x"00",x"00"),
  1972 => (x"66",x"7f",x"19",x"09"),
  1973 => (x"6f",x"26",x"00",x"00"),
  1974 => (x"32",x"7b",x"59",x"4d"),
  1975 => (x"01",x"01",x"00",x"00"),
  1976 => (x"01",x"01",x"7f",x"7f"),
  1977 => (x"7f",x"3f",x"00",x"00"),
  1978 => (x"3f",x"7f",x"40",x"40"),
  1979 => (x"3f",x"0f",x"00",x"00"),
  1980 => (x"0f",x"3f",x"70",x"70"),
  1981 => (x"30",x"7f",x"7f",x"00"),
  1982 => (x"7f",x"7f",x"30",x"18"),
  1983 => (x"36",x"63",x"41",x"00"),
  1984 => (x"63",x"36",x"1c",x"1c"),
  1985 => (x"06",x"03",x"01",x"41"),
  1986 => (x"03",x"06",x"7c",x"7c"),
  1987 => (x"59",x"71",x"61",x"01"),
  1988 => (x"41",x"43",x"47",x"4d"),
  1989 => (x"7f",x"00",x"00",x"00"),
  1990 => (x"00",x"41",x"41",x"7f"),
  1991 => (x"06",x"03",x"01",x"00"),
  1992 => (x"60",x"30",x"18",x"0c"),
  1993 => (x"41",x"00",x"00",x"40"),
  1994 => (x"00",x"7f",x"7f",x"41"),
  1995 => (x"06",x"0c",x"08",x"00"),
  1996 => (x"08",x"0c",x"06",x"03"),
  1997 => (x"80",x"80",x"80",x"00"),
  1998 => (x"80",x"80",x"80",x"80"),
  1999 => (x"00",x"00",x"00",x"00"),
  2000 => (x"00",x"04",x"07",x"03"),
  2001 => (x"74",x"20",x"00",x"00"),
  2002 => (x"78",x"7c",x"54",x"54"),
  2003 => (x"7f",x"7f",x"00",x"00"),
  2004 => (x"38",x"7c",x"44",x"44"),
  2005 => (x"7c",x"38",x"00",x"00"),
  2006 => (x"00",x"44",x"44",x"44"),
  2007 => (x"7c",x"38",x"00",x"00"),
  2008 => (x"7f",x"7f",x"44",x"44"),
  2009 => (x"7c",x"38",x"00",x"00"),
  2010 => (x"18",x"5c",x"54",x"54"),
  2011 => (x"7e",x"04",x"00",x"00"),
  2012 => (x"00",x"05",x"05",x"7f"),
  2013 => (x"bc",x"18",x"00",x"00"),
  2014 => (x"7c",x"fc",x"a4",x"a4"),
  2015 => (x"7f",x"7f",x"00",x"00"),
  2016 => (x"78",x"7c",x"04",x"04"),
  2017 => (x"00",x"00",x"00",x"00"),
  2018 => (x"00",x"40",x"7d",x"3d"),
  2019 => (x"80",x"80",x"00",x"00"),
  2020 => (x"00",x"7d",x"fd",x"80"),
  2021 => (x"7f",x"7f",x"00",x"00"),
  2022 => (x"44",x"6c",x"38",x"10"),
  2023 => (x"00",x"00",x"00",x"00"),
  2024 => (x"00",x"40",x"7f",x"3f"),
  2025 => (x"0c",x"7c",x"7c",x"00"),
  2026 => (x"78",x"7c",x"0c",x"18"),
  2027 => (x"7c",x"7c",x"00",x"00"),
  2028 => (x"78",x"7c",x"04",x"04"),
  2029 => (x"7c",x"38",x"00",x"00"),
  2030 => (x"38",x"7c",x"44",x"44"),
  2031 => (x"fc",x"fc",x"00",x"00"),
  2032 => (x"18",x"3c",x"24",x"24"),
  2033 => (x"3c",x"18",x"00",x"00"),
  2034 => (x"fc",x"fc",x"24",x"24"),
  2035 => (x"7c",x"7c",x"00",x"00"),
  2036 => (x"08",x"0c",x"04",x"04"),
  2037 => (x"5c",x"48",x"00",x"00"),
  2038 => (x"20",x"74",x"54",x"54"),
  2039 => (x"3f",x"04",x"00",x"00"),
  2040 => (x"00",x"44",x"44",x"7f"),
  2041 => (x"7c",x"3c",x"00",x"00"),
  2042 => (x"7c",x"7c",x"40",x"40"),
  2043 => (x"3c",x"1c",x"00",x"00"),
  2044 => (x"1c",x"3c",x"60",x"60"),
  2045 => (x"60",x"7c",x"3c",x"00"),
  2046 => (x"3c",x"7c",x"60",x"30"),
  2047 => (x"38",x"6c",x"44",x"00"),
  2048 => (x"44",x"6c",x"38",x"10"),
  2049 => (x"bc",x"1c",x"00",x"00"),
  2050 => (x"1c",x"3c",x"60",x"e0"),
  2051 => (x"64",x"44",x"00",x"00"),
  2052 => (x"44",x"4c",x"5c",x"74"),
  2053 => (x"08",x"08",x"00",x"00"),
  2054 => (x"41",x"41",x"77",x"3e"),
  2055 => (x"00",x"00",x"00",x"00"),
  2056 => (x"00",x"00",x"7f",x"7f"),
  2057 => (x"41",x"41",x"00",x"00"),
  2058 => (x"08",x"08",x"3e",x"77"),
  2059 => (x"01",x"01",x"02",x"00"),
  2060 => (x"01",x"02",x"02",x"03"),
  2061 => (x"7f",x"7f",x"7f",x"00"),
  2062 => (x"7f",x"7f",x"7f",x"7f"),
  2063 => (x"1c",x"08",x"08",x"00"),
  2064 => (x"7f",x"3e",x"3e",x"1c"),
  2065 => (x"3e",x"7f",x"7f",x"7f"),
  2066 => (x"08",x"1c",x"1c",x"3e"),
  2067 => (x"18",x"10",x"00",x"08"),
  2068 => (x"10",x"18",x"7c",x"7c"),
  2069 => (x"30",x"10",x"00",x"00"),
  2070 => (x"10",x"30",x"7c",x"7c"),
  2071 => (x"60",x"30",x"10",x"00"),
  2072 => (x"06",x"1e",x"78",x"60"),
  2073 => (x"3c",x"66",x"42",x"00"),
  2074 => (x"42",x"66",x"3c",x"18"),
  2075 => (x"6a",x"38",x"78",x"00"),
  2076 => (x"38",x"6c",x"c6",x"c2"),
  2077 => (x"00",x"00",x"60",x"00"),
  2078 => (x"60",x"00",x"00",x"60"),
  2079 => (x"5b",x"5e",x"0e",x"00"),
  2080 => (x"1e",x"0e",x"5d",x"5c"),
  2081 => (x"eb",x"c2",x"4c",x"71"),
  2082 => (x"c0",x"4d",x"bf",x"d6"),
  2083 => (x"74",x"1e",x"c0",x"4b"),
  2084 => (x"87",x"c7",x"02",x"ab"),
  2085 => (x"c0",x"48",x"a6",x"c4"),
  2086 => (x"c4",x"87",x"c5",x"78"),
  2087 => (x"78",x"c1",x"48",x"a6"),
  2088 => (x"73",x"1e",x"66",x"c4"),
  2089 => (x"87",x"df",x"ee",x"49"),
  2090 => (x"e0",x"c0",x"86",x"c8"),
  2091 => (x"87",x"ef",x"ef",x"49"),
  2092 => (x"6a",x"4a",x"a5",x"c4"),
  2093 => (x"87",x"f0",x"f0",x"49"),
  2094 => (x"cb",x"87",x"c6",x"f1"),
  2095 => (x"c8",x"83",x"c1",x"85"),
  2096 => (x"ff",x"04",x"ab",x"b7"),
  2097 => (x"26",x"26",x"87",x"c7"),
  2098 => (x"26",x"4c",x"26",x"4d"),
  2099 => (x"1e",x"4f",x"26",x"4b"),
  2100 => (x"eb",x"c2",x"4a",x"71"),
  2101 => (x"eb",x"c2",x"5a",x"da"),
  2102 => (x"78",x"c7",x"48",x"da"),
  2103 => (x"87",x"dd",x"fe",x"49"),
  2104 => (x"73",x"1e",x"4f",x"26"),
  2105 => (x"c0",x"4a",x"71",x"1e"),
  2106 => (x"d3",x"03",x"aa",x"b7"),
  2107 => (x"f2",x"d0",x"c2",x"87"),
  2108 => (x"87",x"c4",x"05",x"bf"),
  2109 => (x"87",x"c2",x"4b",x"c1"),
  2110 => (x"d0",x"c2",x"4b",x"c0"),
  2111 => (x"87",x"c4",x"5b",x"f6"),
  2112 => (x"5a",x"f6",x"d0",x"c2"),
  2113 => (x"bf",x"f2",x"d0",x"c2"),
  2114 => (x"c1",x"9a",x"c1",x"4a"),
  2115 => (x"ec",x"49",x"a2",x"c0"),
  2116 => (x"48",x"fc",x"87",x"e8"),
  2117 => (x"bf",x"f2",x"d0",x"c2"),
  2118 => (x"87",x"ef",x"fe",x"78"),
  2119 => (x"c4",x"4a",x"71",x"1e"),
  2120 => (x"49",x"72",x"1e",x"66"),
  2121 => (x"26",x"87",x"f5",x"e9"),
  2122 => (x"c2",x"1e",x"4f",x"26"),
  2123 => (x"49",x"bf",x"f2",x"d0"),
  2124 => (x"c2",x"87",x"f3",x"e6"),
  2125 => (x"e8",x"48",x"ce",x"eb"),
  2126 => (x"eb",x"c2",x"78",x"bf"),
  2127 => (x"bf",x"ec",x"48",x"ca"),
  2128 => (x"ce",x"eb",x"c2",x"78"),
  2129 => (x"c3",x"49",x"4a",x"bf"),
  2130 => (x"b7",x"c8",x"99",x"ff"),
  2131 => (x"71",x"48",x"72",x"2a"),
  2132 => (x"d6",x"eb",x"c2",x"b0"),
  2133 => (x"0e",x"4f",x"26",x"58"),
  2134 => (x"5d",x"5c",x"5b",x"5e"),
  2135 => (x"ff",x"4b",x"71",x"0e"),
  2136 => (x"eb",x"c2",x"87",x"c8"),
  2137 => (x"50",x"c0",x"48",x"c9"),
  2138 => (x"d9",x"e6",x"49",x"73"),
  2139 => (x"4c",x"49",x"70",x"87"),
  2140 => (x"ee",x"cb",x"9c",x"c2"),
  2141 => (x"87",x"c2",x"cb",x"49"),
  2142 => (x"c2",x"4d",x"49",x"70"),
  2143 => (x"bf",x"97",x"c9",x"eb"),
  2144 => (x"87",x"e2",x"c1",x"05"),
  2145 => (x"c2",x"49",x"66",x"d0"),
  2146 => (x"99",x"bf",x"d2",x"eb"),
  2147 => (x"d4",x"87",x"d6",x"05"),
  2148 => (x"eb",x"c2",x"49",x"66"),
  2149 => (x"05",x"99",x"bf",x"ca"),
  2150 => (x"49",x"73",x"87",x"cb"),
  2151 => (x"70",x"87",x"e7",x"e5"),
  2152 => (x"c1",x"c1",x"02",x"98"),
  2153 => (x"fe",x"4c",x"c1",x"87"),
  2154 => (x"49",x"75",x"87",x"c0"),
  2155 => (x"70",x"87",x"d7",x"ca"),
  2156 => (x"87",x"c6",x"02",x"98"),
  2157 => (x"48",x"c9",x"eb",x"c2"),
  2158 => (x"eb",x"c2",x"50",x"c1"),
  2159 => (x"05",x"bf",x"97",x"c9"),
  2160 => (x"c2",x"87",x"e3",x"c0"),
  2161 => (x"49",x"bf",x"d2",x"eb"),
  2162 => (x"05",x"99",x"66",x"d0"),
  2163 => (x"c2",x"87",x"d6",x"ff"),
  2164 => (x"49",x"bf",x"ca",x"eb"),
  2165 => (x"05",x"99",x"66",x"d4"),
  2166 => (x"73",x"87",x"ca",x"ff"),
  2167 => (x"87",x"e6",x"e4",x"49"),
  2168 => (x"fe",x"05",x"98",x"70"),
  2169 => (x"48",x"74",x"87",x"ff"),
  2170 => (x"0e",x"87",x"dc",x"fb"),
  2171 => (x"5d",x"5c",x"5b",x"5e"),
  2172 => (x"c0",x"86",x"f4",x"0e"),
  2173 => (x"bf",x"ec",x"4c",x"4d"),
  2174 => (x"48",x"a6",x"c4",x"7e"),
  2175 => (x"bf",x"d6",x"eb",x"c2"),
  2176 => (x"c0",x"1e",x"c1",x"78"),
  2177 => (x"fd",x"49",x"c7",x"1e"),
  2178 => (x"86",x"c8",x"87",x"cd"),
  2179 => (x"cd",x"02",x"98",x"70"),
  2180 => (x"fb",x"49",x"ff",x"87"),
  2181 => (x"da",x"c1",x"87",x"cc"),
  2182 => (x"87",x"ea",x"e3",x"49"),
  2183 => (x"eb",x"c2",x"4d",x"c1"),
  2184 => (x"02",x"bf",x"97",x"c9"),
  2185 => (x"d2",x"cd",x"87",x"c3"),
  2186 => (x"ce",x"eb",x"c2",x"87"),
  2187 => (x"d0",x"c2",x"4b",x"bf"),
  2188 => (x"c0",x"05",x"bf",x"f2"),
  2189 => (x"fd",x"c3",x"87",x"e9"),
  2190 => (x"87",x"ca",x"e3",x"49"),
  2191 => (x"e3",x"49",x"fa",x"c3"),
  2192 => (x"49",x"73",x"87",x"c4"),
  2193 => (x"71",x"99",x"ff",x"c3"),
  2194 => (x"fb",x"49",x"c0",x"1e"),
  2195 => (x"49",x"73",x"87",x"ce"),
  2196 => (x"71",x"29",x"b7",x"c8"),
  2197 => (x"fb",x"49",x"c1",x"1e"),
  2198 => (x"86",x"c8",x"87",x"c2"),
  2199 => (x"c2",x"87",x"f9",x"c5"),
  2200 => (x"4b",x"bf",x"d2",x"eb"),
  2201 => (x"87",x"dd",x"02",x"9b"),
  2202 => (x"bf",x"ee",x"d0",x"c2"),
  2203 => (x"87",x"d6",x"c7",x"49"),
  2204 => (x"c4",x"05",x"98",x"70"),
  2205 => (x"d2",x"4b",x"c0",x"87"),
  2206 => (x"49",x"e0",x"c2",x"87"),
  2207 => (x"c2",x"87",x"fb",x"c6"),
  2208 => (x"c6",x"58",x"f2",x"d0"),
  2209 => (x"ee",x"d0",x"c2",x"87"),
  2210 => (x"73",x"78",x"c0",x"48"),
  2211 => (x"05",x"99",x"c2",x"49"),
  2212 => (x"eb",x"c3",x"87",x"cd"),
  2213 => (x"87",x"ee",x"e1",x"49"),
  2214 => (x"99",x"c2",x"49",x"70"),
  2215 => (x"fb",x"87",x"c2",x"02"),
  2216 => (x"c1",x"49",x"73",x"4c"),
  2217 => (x"87",x"cd",x"05",x"99"),
  2218 => (x"e1",x"49",x"f4",x"c3"),
  2219 => (x"49",x"70",x"87",x"d8"),
  2220 => (x"c2",x"02",x"99",x"c2"),
  2221 => (x"73",x"4c",x"fa",x"87"),
  2222 => (x"05",x"99",x"c8",x"49"),
  2223 => (x"f5",x"c3",x"87",x"cd"),
  2224 => (x"87",x"c2",x"e1",x"49"),
  2225 => (x"99",x"c2",x"49",x"70"),
  2226 => (x"c2",x"87",x"d4",x"02"),
  2227 => (x"02",x"bf",x"da",x"eb"),
  2228 => (x"c1",x"48",x"87",x"c9"),
  2229 => (x"de",x"eb",x"c2",x"88"),
  2230 => (x"ff",x"87",x"c2",x"58"),
  2231 => (x"73",x"4d",x"c1",x"4c"),
  2232 => (x"05",x"99",x"c4",x"49"),
  2233 => (x"f2",x"c3",x"87",x"cd"),
  2234 => (x"87",x"da",x"e0",x"49"),
  2235 => (x"99",x"c2",x"49",x"70"),
  2236 => (x"c2",x"87",x"db",x"02"),
  2237 => (x"7e",x"bf",x"da",x"eb"),
  2238 => (x"a8",x"b7",x"c7",x"48"),
  2239 => (x"6e",x"87",x"cb",x"03"),
  2240 => (x"c2",x"80",x"c1",x"48"),
  2241 => (x"c0",x"58",x"de",x"eb"),
  2242 => (x"4c",x"fe",x"87",x"c2"),
  2243 => (x"fd",x"c3",x"4d",x"c1"),
  2244 => (x"f1",x"df",x"ff",x"49"),
  2245 => (x"c2",x"49",x"70",x"87"),
  2246 => (x"87",x"d5",x"02",x"99"),
  2247 => (x"bf",x"da",x"eb",x"c2"),
  2248 => (x"87",x"c9",x"c0",x"02"),
  2249 => (x"48",x"da",x"eb",x"c2"),
  2250 => (x"c2",x"c0",x"78",x"c0"),
  2251 => (x"c1",x"4c",x"fd",x"87"),
  2252 => (x"49",x"fa",x"c3",x"4d"),
  2253 => (x"87",x"ce",x"df",x"ff"),
  2254 => (x"99",x"c2",x"49",x"70"),
  2255 => (x"c2",x"87",x"d9",x"02"),
  2256 => (x"48",x"bf",x"da",x"eb"),
  2257 => (x"03",x"a8",x"b7",x"c7"),
  2258 => (x"c2",x"87",x"c9",x"c0"),
  2259 => (x"c7",x"48",x"da",x"eb"),
  2260 => (x"87",x"c2",x"c0",x"78"),
  2261 => (x"4d",x"c1",x"4c",x"fc"),
  2262 => (x"03",x"ac",x"b7",x"c0"),
  2263 => (x"c4",x"87",x"d1",x"c0"),
  2264 => (x"d8",x"c1",x"4a",x"66"),
  2265 => (x"c0",x"02",x"6a",x"82"),
  2266 => (x"4b",x"6a",x"87",x"c6"),
  2267 => (x"0f",x"73",x"49",x"74"),
  2268 => (x"f0",x"c3",x"1e",x"c0"),
  2269 => (x"49",x"da",x"c1",x"1e"),
  2270 => (x"c8",x"87",x"dc",x"f7"),
  2271 => (x"02",x"98",x"70",x"86"),
  2272 => (x"c8",x"87",x"e2",x"c0"),
  2273 => (x"eb",x"c2",x"48",x"a6"),
  2274 => (x"c8",x"78",x"bf",x"da"),
  2275 => (x"91",x"cb",x"49",x"66"),
  2276 => (x"71",x"48",x"66",x"c4"),
  2277 => (x"6e",x"7e",x"70",x"80"),
  2278 => (x"c8",x"c0",x"02",x"bf"),
  2279 => (x"4b",x"bf",x"6e",x"87"),
  2280 => (x"73",x"49",x"66",x"c8"),
  2281 => (x"02",x"9d",x"75",x"0f"),
  2282 => (x"c2",x"87",x"c8",x"c0"),
  2283 => (x"49",x"bf",x"da",x"eb"),
  2284 => (x"c2",x"87",x"ca",x"f3"),
  2285 => (x"02",x"bf",x"f6",x"d0"),
  2286 => (x"49",x"87",x"dd",x"c0"),
  2287 => (x"70",x"87",x"c7",x"c2"),
  2288 => (x"d3",x"c0",x"02",x"98"),
  2289 => (x"da",x"eb",x"c2",x"87"),
  2290 => (x"f0",x"f2",x"49",x"bf"),
  2291 => (x"f4",x"49",x"c0",x"87"),
  2292 => (x"d0",x"c2",x"87",x"d0"),
  2293 => (x"78",x"c0",x"48",x"f6"),
  2294 => (x"ea",x"f3",x"8e",x"f4"),
  2295 => (x"5b",x"5e",x"0e",x"87"),
  2296 => (x"1e",x"0e",x"5d",x"5c"),
  2297 => (x"eb",x"c2",x"4c",x"71"),
  2298 => (x"c1",x"49",x"bf",x"d6"),
  2299 => (x"c1",x"4d",x"a1",x"cd"),
  2300 => (x"7e",x"69",x"81",x"d1"),
  2301 => (x"cf",x"02",x"9c",x"74"),
  2302 => (x"4b",x"a5",x"c4",x"87"),
  2303 => (x"eb",x"c2",x"7b",x"74"),
  2304 => (x"f3",x"49",x"bf",x"d6"),
  2305 => (x"7b",x"6e",x"87",x"c9"),
  2306 => (x"c4",x"05",x"9c",x"74"),
  2307 => (x"c2",x"4b",x"c0",x"87"),
  2308 => (x"73",x"4b",x"c1",x"87"),
  2309 => (x"87",x"ca",x"f3",x"49"),
  2310 => (x"c7",x"02",x"66",x"d4"),
  2311 => (x"87",x"da",x"49",x"87"),
  2312 => (x"87",x"c2",x"4a",x"70"),
  2313 => (x"d0",x"c2",x"4a",x"c0"),
  2314 => (x"f2",x"26",x"5a",x"fa"),
  2315 => (x"00",x"00",x"87",x"d9"),
  2316 => (x"00",x"00",x"00",x"00"),
  2317 => (x"00",x"00",x"00",x"00"),
  2318 => (x"71",x"1e",x"00",x"00"),
  2319 => (x"bf",x"c8",x"ff",x"4a"),
  2320 => (x"48",x"a1",x"72",x"49"),
  2321 => (x"ff",x"1e",x"4f",x"26"),
  2322 => (x"fe",x"89",x"bf",x"c8"),
  2323 => (x"c0",x"c0",x"c0",x"c0"),
  2324 => (x"c4",x"01",x"a9",x"c0"),
  2325 => (x"c2",x"4a",x"c0",x"87"),
  2326 => (x"72",x"4a",x"c1",x"87"),
  2327 => (x"0e",x"4f",x"26",x"48"),
  2328 => (x"5d",x"5c",x"5b",x"5e"),
  2329 => (x"7e",x"71",x"1e",x"0e"),
  2330 => (x"6e",x"4b",x"d4",x"ff"),
  2331 => (x"de",x"eb",x"c2",x"1e"),
  2332 => (x"d8",x"cf",x"fe",x"49"),
  2333 => (x"70",x"86",x"c4",x"87"),
  2334 => (x"c3",x"02",x"9d",x"4d"),
  2335 => (x"eb",x"c2",x"87",x"c3"),
  2336 => (x"6e",x"4c",x"bf",x"e6"),
  2337 => (x"d0",x"e2",x"fe",x"49"),
  2338 => (x"48",x"d0",x"ff",x"87"),
  2339 => (x"c1",x"78",x"c5",x"c8"),
  2340 => (x"4a",x"c0",x"7b",x"d6"),
  2341 => (x"82",x"c1",x"7b",x"15"),
  2342 => (x"aa",x"b7",x"e0",x"c0"),
  2343 => (x"ff",x"87",x"f5",x"04"),
  2344 => (x"78",x"c4",x"48",x"d0"),
  2345 => (x"c1",x"78",x"c5",x"c8"),
  2346 => (x"7b",x"c1",x"7b",x"d3"),
  2347 => (x"9c",x"74",x"78",x"c4"),
  2348 => (x"87",x"fc",x"c1",x"02"),
  2349 => (x"7e",x"ce",x"da",x"c2"),
  2350 => (x"8c",x"4d",x"c0",x"c8"),
  2351 => (x"03",x"ac",x"b7",x"c0"),
  2352 => (x"c0",x"c8",x"87",x"c6"),
  2353 => (x"4c",x"c0",x"4d",x"a4"),
  2354 => (x"97",x"ff",x"e6",x"c2"),
  2355 => (x"99",x"d0",x"49",x"bf"),
  2356 => (x"c0",x"87",x"d2",x"02"),
  2357 => (x"de",x"eb",x"c2",x"1e"),
  2358 => (x"cc",x"d1",x"fe",x"49"),
  2359 => (x"70",x"86",x"c4",x"87"),
  2360 => (x"ef",x"c0",x"4a",x"49"),
  2361 => (x"ce",x"da",x"c2",x"87"),
  2362 => (x"de",x"eb",x"c2",x"1e"),
  2363 => (x"f8",x"d0",x"fe",x"49"),
  2364 => (x"70",x"86",x"c4",x"87"),
  2365 => (x"d0",x"ff",x"4a",x"49"),
  2366 => (x"78",x"c5",x"c8",x"48"),
  2367 => (x"6e",x"7b",x"d4",x"c1"),
  2368 => (x"6e",x"7b",x"bf",x"97"),
  2369 => (x"70",x"80",x"c1",x"48"),
  2370 => (x"05",x"8d",x"c1",x"7e"),
  2371 => (x"ff",x"87",x"f0",x"ff"),
  2372 => (x"78",x"c4",x"48",x"d0"),
  2373 => (x"c5",x"05",x"9a",x"72"),
  2374 => (x"c0",x"48",x"c0",x"87"),
  2375 => (x"1e",x"c1",x"87",x"e5"),
  2376 => (x"49",x"de",x"eb",x"c2"),
  2377 => (x"87",x"e0",x"ce",x"fe"),
  2378 => (x"9c",x"74",x"86",x"c4"),
  2379 => (x"87",x"c4",x"fe",x"05"),
  2380 => (x"c8",x"48",x"d0",x"ff"),
  2381 => (x"d3",x"c1",x"78",x"c5"),
  2382 => (x"c4",x"7b",x"c0",x"7b"),
  2383 => (x"c2",x"48",x"c1",x"78"),
  2384 => (x"26",x"48",x"c0",x"87"),
  2385 => (x"4c",x"26",x"4d",x"26"),
  2386 => (x"4f",x"26",x"4b",x"26"),
  2387 => (x"71",x"1e",x"73",x"1e"),
  2388 => (x"02",x"66",x"c8",x"4a"),
  2389 => (x"c1",x"4b",x"87",x"ce"),
  2390 => (x"ce",x"02",x"8b",x"d3"),
  2391 => (x"02",x"8b",x"c1",x"87"),
  2392 => (x"87",x"d3",x"87",x"d0"),
  2393 => (x"f6",x"fb",x"49",x"72"),
  2394 => (x"72",x"87",x"cc",x"87"),
  2395 => (x"87",x"ca",x"c2",x"49"),
  2396 => (x"49",x"72",x"87",x"c5"),
  2397 => (x"ff",x"87",x"f6",x"c2"),
  2398 => (x"1e",x"00",x"87",x"ce"),
  2399 => (x"bf",x"e2",x"d9",x"c2"),
  2400 => (x"c2",x"b9",x"c1",x"49"),
  2401 => (x"ff",x"59",x"e6",x"d9"),
  2402 => (x"ff",x"c3",x"48",x"d4"),
  2403 => (x"48",x"d0",x"ff",x"78"),
  2404 => (x"ff",x"78",x"e1",x"c8"),
  2405 => (x"78",x"c1",x"48",x"d4"),
  2406 => (x"78",x"71",x"31",x"c4"),
  2407 => (x"c0",x"48",x"d0",x"ff"),
  2408 => (x"4f",x"26",x"78",x"e0"),
  2409 => (x"fd",x"d6",x"c2",x"1e"),
  2410 => (x"de",x"eb",x"c2",x"1e"),
  2411 => (x"dc",x"ca",x"fe",x"49"),
  2412 => (x"70",x"86",x"c4",x"87"),
  2413 => (x"87",x"c3",x"02",x"98"),
  2414 => (x"26",x"87",x"c0",x"ff"),
  2415 => (x"4b",x"35",x"31",x"4f"),
  2416 => (x"20",x"20",x"5a",x"48"),
  2417 => (x"47",x"46",x"43",x"20"),
  2418 => (x"4a",x"71",x"1e",x"00"),
  2419 => (x"c2",x"49",x"a2",x"c4"),
  2420 => (x"6a",x"48",x"f5",x"ea"),
  2421 => (x"c1",x"49",x"69",x"78"),
  2422 => (x"e6",x"d9",x"c2",x"b9"),
  2423 => (x"87",x"db",x"fe",x"59"),
  2424 => (x"87",x"d9",x"d7",x"ff"),
  2425 => (x"4f",x"26",x"48",x"c1"),
  2426 => (x"c4",x"4a",x"71",x"1e"),
  2427 => (x"ea",x"c2",x"49",x"a2"),
  2428 => (x"c2",x"7a",x"bf",x"f5"),
  2429 => (x"79",x"bf",x"e2",x"d9"),
  2430 => (x"71",x"1e",x"4f",x"26"),
  2431 => (x"eb",x"c2",x"1e",x"4a"),
  2432 => (x"c9",x"fe",x"49",x"de"),
  2433 => (x"86",x"c4",x"87",x"c7"),
  2434 => (x"dc",x"02",x"98",x"70"),
  2435 => (x"ce",x"da",x"c2",x"87"),
  2436 => (x"de",x"eb",x"c2",x"1e"),
  2437 => (x"d0",x"cc",x"fe",x"49"),
  2438 => (x"70",x"86",x"c4",x"87"),
  2439 => (x"87",x"c9",x"02",x"98"),
  2440 => (x"49",x"ce",x"da",x"c2"),
  2441 => (x"c2",x"87",x"e2",x"fe"),
  2442 => (x"26",x"48",x"c0",x"87"),
  2443 => (x"4a",x"71",x"1e",x"4f"),
  2444 => (x"de",x"eb",x"c2",x"1e"),
  2445 => (x"d4",x"c8",x"fe",x"49"),
  2446 => (x"70",x"86",x"c4",x"87"),
  2447 => (x"87",x"de",x"02",x"98"),
  2448 => (x"49",x"ce",x"da",x"c2"),
  2449 => (x"c2",x"87",x"e1",x"fe"),
  2450 => (x"c2",x"1e",x"ce",x"da"),
  2451 => (x"fe",x"49",x"de",x"eb"),
  2452 => (x"c4",x"87",x"d9",x"cc"),
  2453 => (x"02",x"98",x"70",x"86"),
  2454 => (x"48",x"c1",x"87",x"c4"),
  2455 => (x"48",x"c0",x"87",x"c2"),
  2456 => (x"00",x"00",x"4f",x"26"),
  2457 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

