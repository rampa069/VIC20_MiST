library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f4ebc287",
    12 => x"86c0c64e",
    13 => x"49f4ebc2",
    14 => x"48e8d9c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e0de",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48111e4f",
    50 => x"7808d4ff",
    51 => x"c14866c4",
    52 => x"58a6c888",
    53 => x"ed059870",
    54 => x"1e4f2687",
    55 => x"c348d4ff",
    56 => x"516878ff",
    57 => x"c14866c4",
    58 => x"58a6c888",
    59 => x"eb059870",
    60 => x"1e4f2687",
    61 => x"d4ff1e73",
    62 => x"7bffc34b",
    63 => x"ffc34a6b",
    64 => x"c8496b7b",
    65 => x"c3b17232",
    66 => x"4a6b7bff",
    67 => x"b27131c8",
    68 => x"6b7bffc3",
    69 => x"7232c849",
    70 => x"c44871b1",
    71 => x"264d2687",
    72 => x"264b264c",
    73 => x"5b5e0e4f",
    74 => x"710e5d5c",
    75 => x"4cd4ff4a",
    76 => x"ffc34972",
    77 => x"c27c7199",
    78 => x"05bfe8d9",
    79 => x"66d087c8",
    80 => x"d430c948",
    81 => x"66d058a6",
    82 => x"c329d849",
    83 => x"7c7199ff",
    84 => x"d04966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"c329c849",
    88 => x"7c7199ff",
    89 => x"c34966d0",
    90 => x"7c7199ff",
    91 => x"29d04972",
    92 => x"7199ffc3",
    93 => x"c94b6c7c",
    94 => x"c34dfff0",
    95 => x"d005abff",
    96 => x"7cffc387",
    97 => x"8dc14b6c",
    98 => x"c387c602",
    99 => x"f002abff",
   100 => x"fe487387",
   101 => x"c01e87c7",
   102 => x"48d4ff49",
   103 => x"c178ffc3",
   104 => x"b7c8c381",
   105 => x"87f104a9",
   106 => x"731e4f26",
   107 => x"c487e71e",
   108 => x"c04bdff8",
   109 => x"f0ffc01e",
   110 => x"fd49f7c1",
   111 => x"86c487e7",
   112 => x"c005a8c1",
   113 => x"d4ff87ea",
   114 => x"78ffc348",
   115 => x"c0c0c0c1",
   116 => x"c01ec0c0",
   117 => x"e9c1f0e1",
   118 => x"87c9fd49",
   119 => x"987086c4",
   120 => x"ff87ca05",
   121 => x"ffc348d4",
   122 => x"cb48c178",
   123 => x"87e6fe87",
   124 => x"fe058bc1",
   125 => x"48c087fd",
   126 => x"1e87e6fc",
   127 => x"d4ff1e73",
   128 => x"78ffc348",
   129 => x"1ec04bd3",
   130 => x"c1f0ffc0",
   131 => x"d4fc49c1",
   132 => x"7086c487",
   133 => x"87ca0598",
   134 => x"c348d4ff",
   135 => x"48c178ff",
   136 => x"f1fd87cb",
   137 => x"058bc187",
   138 => x"c087dbff",
   139 => x"87f1fb48",
   140 => x"5c5b5e0e",
   141 => x"4cd4ff0e",
   142 => x"c687dbfd",
   143 => x"e1c01eea",
   144 => x"49c8c1f0",
   145 => x"c487defb",
   146 => x"02a8c186",
   147 => x"eafe87c8",
   148 => x"c148c087",
   149 => x"dafa87e2",
   150 => x"cf497087",
   151 => x"c699ffff",
   152 => x"c802a9ea",
   153 => x"87d3fe87",
   154 => x"cbc148c0",
   155 => x"7cffc387",
   156 => x"fc4bf1c0",
   157 => x"987087f4",
   158 => x"87ebc002",
   159 => x"ffc01ec0",
   160 => x"49fac1f0",
   161 => x"c487defa",
   162 => x"05987086",
   163 => x"ffc387d9",
   164 => x"c3496c7c",
   165 => x"7c7c7cff",
   166 => x"99c0c17c",
   167 => x"c187c402",
   168 => x"c087d548",
   169 => x"c287d148",
   170 => x"87c405ab",
   171 => x"87c848c0",
   172 => x"fe058bc1",
   173 => x"48c087fd",
   174 => x"1e87e4f9",
   175 => x"d9c21e73",
   176 => x"78c148e8",
   177 => x"d0ff4bc7",
   178 => x"fb78c248",
   179 => x"d0ff87c8",
   180 => x"c078c348",
   181 => x"d0e5c01e",
   182 => x"f949c0c1",
   183 => x"86c487c7",
   184 => x"c105a8c1",
   185 => x"abc24b87",
   186 => x"c087c505",
   187 => x"87f9c048",
   188 => x"ff058bc1",
   189 => x"f7fc87d0",
   190 => x"ecd9c287",
   191 => x"05987058",
   192 => x"1ec187cd",
   193 => x"c1f0ffc0",
   194 => x"d8f849d0",
   195 => x"ff86c487",
   196 => x"ffc348d4",
   197 => x"87e0c478",
   198 => x"58f0d9c2",
   199 => x"c248d0ff",
   200 => x"48d4ff78",
   201 => x"c178ffc3",
   202 => x"87f5f748",
   203 => x"5c5b5e0e",
   204 => x"4a710e5d",
   205 => x"ff4dffc3",
   206 => x"7c754cd4",
   207 => x"c448d0ff",
   208 => x"7c7578c3",
   209 => x"ffc01e72",
   210 => x"49d8c1f0",
   211 => x"c487d6f7",
   212 => x"02987086",
   213 => x"48c087c5",
   214 => x"7587f0c0",
   215 => x"7cfec37c",
   216 => x"d41ec0c8",
   217 => x"dcf54966",
   218 => x"7586c487",
   219 => x"757c757c",
   220 => x"e0dad87c",
   221 => x"6c7c754b",
   222 => x"c5059949",
   223 => x"058bc187",
   224 => x"7c7587f3",
   225 => x"c248d0ff",
   226 => x"f648c178",
   227 => x"ff1e87cf",
   228 => x"d0ff4ad4",
   229 => x"78d1c448",
   230 => x"c17affc3",
   231 => x"87f80589",
   232 => x"731e4f26",
   233 => x"c54b711e",
   234 => x"4adfcdee",
   235 => x"c348d4ff",
   236 => x"486878ff",
   237 => x"02a8fec3",
   238 => x"8ac187c5",
   239 => x"7287ed05",
   240 => x"87c5059a",
   241 => x"eac048c0",
   242 => x"029b7387",
   243 => x"66c887cc",
   244 => x"f449731e",
   245 => x"86c487c5",
   246 => x"66c887c6",
   247 => x"87eefe49",
   248 => x"c348d4ff",
   249 => x"737878ff",
   250 => x"87c5059b",
   251 => x"d048d0ff",
   252 => x"f448c178",
   253 => x"731e87eb",
   254 => x"c04a711e",
   255 => x"48d4ff4b",
   256 => x"ff78ffc3",
   257 => x"c3c448d0",
   258 => x"48d4ff78",
   259 => x"7278ffc3",
   260 => x"f0ffc01e",
   261 => x"f449d1c1",
   262 => x"86c487cb",
   263 => x"cd059870",
   264 => x"1ec0c887",
   265 => x"fd4966cc",
   266 => x"86c487f8",
   267 => x"d0ff4b70",
   268 => x"7378c248",
   269 => x"87e9f348",
   270 => x"5c5b5e0e",
   271 => x"1ec00e5d",
   272 => x"c1f0ffc0",
   273 => x"dcf349c9",
   274 => x"c21ed287",
   275 => x"fd49f0d9",
   276 => x"86c887d0",
   277 => x"84c14cc0",
   278 => x"04acb7d2",
   279 => x"d9c287f8",
   280 => x"49bf97f0",
   281 => x"c199c0c3",
   282 => x"c005a9c0",
   283 => x"d9c287e7",
   284 => x"49bf97f7",
   285 => x"d9c231d0",
   286 => x"4abf97f8",
   287 => x"b17232c8",
   288 => x"97f9d9c2",
   289 => x"71b14abf",
   290 => x"ffffcf4c",
   291 => x"84c19cff",
   292 => x"e7c134ca",
   293 => x"f9d9c287",
   294 => x"c149bf97",
   295 => x"c299c631",
   296 => x"bf97fad9",
   297 => x"2ab7c74a",
   298 => x"d9c2b172",
   299 => x"4abf97f5",
   300 => x"c29dcf4d",
   301 => x"bf97f6d9",
   302 => x"ca9ac34a",
   303 => x"f7d9c232",
   304 => x"c24bbf97",
   305 => x"c2b27333",
   306 => x"bf97f8d9",
   307 => x"9bc0c34b",
   308 => x"732bb7c6",
   309 => x"c181c2b2",
   310 => x"70307148",
   311 => x"7548c149",
   312 => x"724d7030",
   313 => x"7184c14c",
   314 => x"b7c0c894",
   315 => x"87cc06ad",
   316 => x"2db734c1",
   317 => x"adb7c0c8",
   318 => x"87f4ff01",
   319 => x"dcf04874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"d6e2c286",
   323 => x"c278c048",
   324 => x"c01eceda",
   325 => x"87defb49",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec948",
   329 => x"7ec14dc0",
   330 => x"bfe4f0c0",
   331 => x"c4dbc249",
   332 => x"4bc8714a",
   333 => x"7087f3ec",
   334 => x"87c20598",
   335 => x"f0c07ec0",
   336 => x"c249bfe0",
   337 => x"714ae0db",
   338 => x"ddec4bc8",
   339 => x"05987087",
   340 => x"7ec087c2",
   341 => x"fdc0026e",
   342 => x"d4e1c287",
   343 => x"e2c24dbf",
   344 => x"7ebf9fcc",
   345 => x"ead6c548",
   346 => x"87c705a8",
   347 => x"bfd4e1c2",
   348 => x"6e87ce4d",
   349 => x"d5e9ca48",
   350 => x"87c502a8",
   351 => x"f1c748c0",
   352 => x"cedac287",
   353 => x"f949751e",
   354 => x"86c487ec",
   355 => x"c5059870",
   356 => x"c748c087",
   357 => x"f0c087dc",
   358 => x"c249bfe0",
   359 => x"714ae0db",
   360 => x"c5eb4bc8",
   361 => x"05987087",
   362 => x"e2c287c8",
   363 => x"78c148d6",
   364 => x"f0c087da",
   365 => x"c249bfe4",
   366 => x"714ac4db",
   367 => x"e9ea4bc8",
   368 => x"02987087",
   369 => x"c087c5c0",
   370 => x"87e6c648",
   371 => x"97cce2c2",
   372 => x"d5c149bf",
   373 => x"cdc005a9",
   374 => x"cde2c287",
   375 => x"c249bf97",
   376 => x"c002a9ea",
   377 => x"48c087c5",
   378 => x"c287c7c6",
   379 => x"bf97ceda",
   380 => x"e9c3487e",
   381 => x"cec002a8",
   382 => x"c3486e87",
   383 => x"c002a8eb",
   384 => x"48c087c5",
   385 => x"c287ebc5",
   386 => x"bf97d9da",
   387 => x"c0059949",
   388 => x"dac287cc",
   389 => x"49bf97da",
   390 => x"c002a9c2",
   391 => x"48c087c5",
   392 => x"c287cfc5",
   393 => x"bf97dbda",
   394 => x"d2e2c248",
   395 => x"484c7058",
   396 => x"e2c288c1",
   397 => x"dac258d6",
   398 => x"49bf97dc",
   399 => x"dac28175",
   400 => x"4abf97dd",
   401 => x"a17232c8",
   402 => x"e3e6c27e",
   403 => x"c2786e48",
   404 => x"bf97deda",
   405 => x"58a6c848",
   406 => x"bfd6e2c2",
   407 => x"87d4c202",
   408 => x"bfe0f0c0",
   409 => x"e0dbc249",
   410 => x"4bc8714a",
   411 => x"7087fbe7",
   412 => x"c5c00298",
   413 => x"c348c087",
   414 => x"e2c287f8",
   415 => x"c24cbfce",
   416 => x"c25cf7e6",
   417 => x"bf97f3da",
   418 => x"c231c849",
   419 => x"bf97f2da",
   420 => x"c249a14a",
   421 => x"bf97f4da",
   422 => x"7232d04a",
   423 => x"dac249a1",
   424 => x"4abf97f5",
   425 => x"a17232d8",
   426 => x"9166c449",
   427 => x"bfe3e6c2",
   428 => x"ebe6c281",
   429 => x"fbdac259",
   430 => x"c84abf97",
   431 => x"fadac232",
   432 => x"a24bbf97",
   433 => x"fcdac24a",
   434 => x"d04bbf97",
   435 => x"4aa27333",
   436 => x"97fddac2",
   437 => x"9bcf4bbf",
   438 => x"a27333d8",
   439 => x"efe6c24a",
   440 => x"ebe6c25a",
   441 => x"8ac24abf",
   442 => x"e6c29274",
   443 => x"a17248ef",
   444 => x"87cac178",
   445 => x"97e0dac2",
   446 => x"31c849bf",
   447 => x"97dfdac2",
   448 => x"49a14abf",
   449 => x"59dee2c2",
   450 => x"bfdae2c2",
   451 => x"c731c549",
   452 => x"29c981ff",
   453 => x"59f7e6c2",
   454 => x"97e5dac2",
   455 => x"32c84abf",
   456 => x"97e4dac2",
   457 => x"4aa24bbf",
   458 => x"6e9266c4",
   459 => x"f3e6c282",
   460 => x"ebe6c25a",
   461 => x"c278c048",
   462 => x"7248e7e6",
   463 => x"e6c278a1",
   464 => x"e6c248f7",
   465 => x"c278bfeb",
   466 => x"c248fbe6",
   467 => x"78bfefe6",
   468 => x"bfd6e2c2",
   469 => x"87c9c002",
   470 => x"30c44874",
   471 => x"c9c07e70",
   472 => x"f3e6c287",
   473 => x"30c448bf",
   474 => x"e2c27e70",
   475 => x"786e48da",
   476 => x"8ef848c1",
   477 => x"4c264d26",
   478 => x"4f264b26",
   479 => x"5c5b5e0e",
   480 => x"4a710e5d",
   481 => x"bfd6e2c2",
   482 => x"7287cb02",
   483 => x"722bc74b",
   484 => x"9cffc14c",
   485 => x"4b7287c9",
   486 => x"4c722bc8",
   487 => x"c29cffc3",
   488 => x"83bfe3e6",
   489 => x"bfdcf0c0",
   490 => x"87d902ab",
   491 => x"5be0f0c0",
   492 => x"1ecedac2",
   493 => x"fdf04973",
   494 => x"7086c487",
   495 => x"87c50598",
   496 => x"e6c048c0",
   497 => x"d6e2c287",
   498 => x"87d202bf",
   499 => x"91c44974",
   500 => x"81cedac2",
   501 => x"ffcf4d69",
   502 => x"9dffffff",
   503 => x"497487cb",
   504 => x"dac291c2",
   505 => x"699f81ce",
   506 => x"fe48754d",
   507 => x"5e0e87c6",
   508 => x"0e5d5c5b",
   509 => x"c04d711e",
   510 => x"c949c11e",
   511 => x"86c487c7",
   512 => x"029c4c70",
   513 => x"c287c0c1",
   514 => x"754adee2",
   515 => x"87ffe049",
   516 => x"c0029870",
   517 => x"4a7487f1",
   518 => x"4bcb4975",
   519 => x"7087e5e1",
   520 => x"e2c00298",
   521 => x"741ec087",
   522 => x"87c7029c",
   523 => x"c048a6c4",
   524 => x"c487c578",
   525 => x"78c148a6",
   526 => x"c84966c4",
   527 => x"86c487c7",
   528 => x"059c4c70",
   529 => x"7487c0ff",
   530 => x"e7fc2648",
   531 => x"5b5e0e87",
   532 => x"1e0e5d5c",
   533 => x"059b4b71",
   534 => x"48c087c5",
   535 => x"c887e5c1",
   536 => x"7dc04da3",
   537 => x"c70266d4",
   538 => x"9766d487",
   539 => x"87c505bf",
   540 => x"cfc148c0",
   541 => x"4966d487",
   542 => x"7087f3fd",
   543 => x"c1029c4c",
   544 => x"a4dc87c0",
   545 => x"da7d6949",
   546 => x"a3c449a4",
   547 => x"7a699f4a",
   548 => x"bfd6e2c2",
   549 => x"d487d202",
   550 => x"699f49a4",
   551 => x"ffffc049",
   552 => x"d0487199",
   553 => x"c27e7030",
   554 => x"6e7ec087",
   555 => x"806a4849",
   556 => x"7bc07a70",
   557 => x"6a49a3cc",
   558 => x"49a3d079",
   559 => x"487479c0",
   560 => x"48c087c2",
   561 => x"87ecfa26",
   562 => x"5c5b5e0e",
   563 => x"4c710e5d",
   564 => x"48dcf0c0",
   565 => x"9c7478ff",
   566 => x"87cac102",
   567 => x"6949a4c8",
   568 => x"87c2c102",
   569 => x"6c4a66d0",
   570 => x"a6d48249",
   571 => x"4d66d05a",
   572 => x"d2e2c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e4c002",
   576 => x"6b4ba4c4",
   577 => x"87f4f949",
   578 => x"e2c27b70",
   579 => x"6c49bfce",
   580 => x"757c7181",
   581 => x"d2e2c2b9",
   582 => x"baff4abf",
   583 => x"99719972",
   584 => x"87dcff05",
   585 => x"cbf97c75",
   586 => x"1e731e87",
   587 => x"029b4b71",
   588 => x"a3c887c7",
   589 => x"c5056949",
   590 => x"c048c087",
   591 => x"e6c287eb",
   592 => x"c44abfe7",
   593 => x"496949a3",
   594 => x"e2c289c2",
   595 => x"7191bfce",
   596 => x"e2c24aa2",
   597 => x"6b49bfd2",
   598 => x"4aa27199",
   599 => x"721e66c8",
   600 => x"87d2ea49",
   601 => x"497086c4",
   602 => x"87ccf848",
   603 => x"711e731e",
   604 => x"c7029b4b",
   605 => x"49a3c887",
   606 => x"87c50569",
   607 => x"ebc048c0",
   608 => x"e7e6c287",
   609 => x"a3c44abf",
   610 => x"c2496949",
   611 => x"cee2c289",
   612 => x"a27191bf",
   613 => x"d2e2c24a",
   614 => x"996b49bf",
   615 => x"c84aa271",
   616 => x"49721e66",
   617 => x"c487c5e6",
   618 => x"48497086",
   619 => x"1e87c9f7",
   620 => x"4b711e73",
   621 => x"e4c0029b",
   622 => x"fbe6c287",
   623 => x"c24a735b",
   624 => x"cee2c28a",
   625 => x"c29249bf",
   626 => x"48bfe7e6",
   627 => x"e6c28072",
   628 => x"487158ff",
   629 => x"e2c230c4",
   630 => x"edc058de",
   631 => x"f7e6c287",
   632 => x"ebe6c248",
   633 => x"e6c278bf",
   634 => x"e6c248fb",
   635 => x"c278bfef",
   636 => x"02bfd6e2",
   637 => x"e2c287c9",
   638 => x"c449bfce",
   639 => x"c287c731",
   640 => x"49bff3e6",
   641 => x"e2c231c4",
   642 => x"ebf559de",
   643 => x"5b5e0e87",
   644 => x"4a710e5c",
   645 => x"9a724bc0",
   646 => x"87e1c002",
   647 => x"9f49a2da",
   648 => x"e2c24b69",
   649 => x"cf02bfd6",
   650 => x"49a2d487",
   651 => x"4c49699f",
   652 => x"9cffffc0",
   653 => x"87c234d0",
   654 => x"49744cc0",
   655 => x"fd4973b3",
   656 => x"f1f487ed",
   657 => x"5b5e0e87",
   658 => x"f40e5d5c",
   659 => x"c04a7186",
   660 => x"029a727e",
   661 => x"dac287d8",
   662 => x"78c048ca",
   663 => x"48c2dac2",
   664 => x"bffbe6c2",
   665 => x"c6dac278",
   666 => x"f7e6c248",
   667 => x"e2c278bf",
   668 => x"50c048eb",
   669 => x"bfdae2c2",
   670 => x"cadac249",
   671 => x"aa714abf",
   672 => x"87ffc303",
   673 => x"99cf4972",
   674 => x"87e0c005",
   675 => x"1ecedac2",
   676 => x"bfc2dac2",
   677 => x"c2dac249",
   678 => x"78a1c148",
   679 => x"87d6e571",
   680 => x"f0c086c4",
   681 => x"dac248d8",
   682 => x"87cc78ce",
   683 => x"bfd8f0c0",
   684 => x"80e0c048",
   685 => x"58dcf0c0",
   686 => x"bfcadac2",
   687 => x"c280c148",
   688 => x"2758ceda",
   689 => x"00000c18",
   690 => x"4dbf97bf",
   691 => x"e2c2029d",
   692 => x"ade5c387",
   693 => x"87dbc202",
   694 => x"bfd8f0c0",
   695 => x"49a3cb4b",
   696 => x"accf4c11",
   697 => x"87d2c105",
   698 => x"99df4975",
   699 => x"91cd89c1",
   700 => x"81dee2c2",
   701 => x"124aa3c1",
   702 => x"4aa3c351",
   703 => x"a3c55112",
   704 => x"c751124a",
   705 => x"51124aa3",
   706 => x"124aa3c9",
   707 => x"4aa3ce51",
   708 => x"a3d05112",
   709 => x"d251124a",
   710 => x"51124aa3",
   711 => x"124aa3d4",
   712 => x"4aa3d651",
   713 => x"a3d85112",
   714 => x"dc51124a",
   715 => x"51124aa3",
   716 => x"124aa3de",
   717 => x"c07ec151",
   718 => x"497487f9",
   719 => x"c00599c8",
   720 => x"497487ea",
   721 => x"d00599d0",
   722 => x"0266dc87",
   723 => x"7387cac0",
   724 => x"0f66dc49",
   725 => x"d3029870",
   726 => x"c0056e87",
   727 => x"e2c287c6",
   728 => x"50c048de",
   729 => x"bfd8f0c0",
   730 => x"87e7c248",
   731 => x"48ebe2c2",
   732 => x"c27e50c0",
   733 => x"49bfdae2",
   734 => x"bfcadac2",
   735 => x"04aa714a",
   736 => x"c287c1fc",
   737 => x"05bffbe6",
   738 => x"c287c8c0",
   739 => x"02bfd6e2",
   740 => x"c087fec1",
   741 => x"ff48dcf0",
   742 => x"c6dac278",
   743 => x"dbef49bf",
   744 => x"c2497087",
   745 => x"c459cada",
   746 => x"dac248a6",
   747 => x"c278bfc6",
   748 => x"02bfd6e2",
   749 => x"c487d8c0",
   750 => x"ffcf4966",
   751 => x"99f8ffff",
   752 => x"c5c002a9",
   753 => x"c04dc087",
   754 => x"4dc187e1",
   755 => x"c487dcc0",
   756 => x"ffcf4966",
   757 => x"02a999f8",
   758 => x"c887c8c0",
   759 => x"78c048a6",
   760 => x"c887c5c0",
   761 => x"78c148a6",
   762 => x"754d66c8",
   763 => x"e0c0059d",
   764 => x"4966c487",
   765 => x"e2c289c2",
   766 => x"914abfce",
   767 => x"bfe7e6c2",
   768 => x"c2dac24a",
   769 => x"78a17248",
   770 => x"48cadac2",
   771 => x"e3f978c0",
   772 => x"f448c087",
   773 => x"87dced8e",
   774 => x"00000000",
   775 => x"ffffffff",
   776 => x"00000c28",
   777 => x"00000c31",
   778 => x"33544146",
   779 => x"20202032",
   780 => x"54414600",
   781 => x"20203631",
   782 => x"ff1e0020",
   783 => x"ffc348d4",
   784 => x"26486878",
   785 => x"d4ff1e4f",
   786 => x"78ffc348",
   787 => x"c848d0ff",
   788 => x"d4ff78e1",
   789 => x"c278d448",
   790 => x"ff48ffe6",
   791 => x"2650bfd4",
   792 => x"d0ff1e4f",
   793 => x"78e0c048",
   794 => x"ff1e4f26",
   795 => x"497087cc",
   796 => x"87c60299",
   797 => x"05a9fbc0",
   798 => x"487187f1",
   799 => x"5e0e4f26",
   800 => x"710e5c5b",
   801 => x"fe4cc04b",
   802 => x"497087f0",
   803 => x"f9c00299",
   804 => x"a9ecc087",
   805 => x"87f2c002",
   806 => x"02a9fbc0",
   807 => x"cc87ebc0",
   808 => x"03acb766",
   809 => x"66d087c7",
   810 => x"7187c202",
   811 => x"02997153",
   812 => x"84c187c2",
   813 => x"7087c3fe",
   814 => x"cd029949",
   815 => x"a9ecc087",
   816 => x"c087c702",
   817 => x"ff05a9fb",
   818 => x"66d087d5",
   819 => x"c087c302",
   820 => x"ecc07b97",
   821 => x"87c405a9",
   822 => x"87c54a74",
   823 => x"0ac04a74",
   824 => x"c248728a",
   825 => x"264d2687",
   826 => x"264b264c",
   827 => x"c9fd1e4f",
   828 => x"c0497087",
   829 => x"04a9b7f0",
   830 => x"f9c087ca",
   831 => x"c301a9b7",
   832 => x"89f0c087",
   833 => x"a9b7c1c1",
   834 => x"c187ca04",
   835 => x"01a9b7da",
   836 => x"f7c087c3",
   837 => x"26487189",
   838 => x"5b5e0e4f",
   839 => x"4a710e5c",
   840 => x"724cd4ff",
   841 => x"87eac049",
   842 => x"029b4b70",
   843 => x"8bc187c2",
   844 => x"c848d0ff",
   845 => x"d5c178c5",
   846 => x"c649737c",
   847 => x"fad5c231",
   848 => x"484abf97",
   849 => x"7c70b071",
   850 => x"c448d0ff",
   851 => x"fe487378",
   852 => x"5e0e87d5",
   853 => x"0e5d5c5b",
   854 => x"4b7186f8",
   855 => x"f8c07ec0",
   856 => x"49bf97f9",
   857 => x"c005a9df",
   858 => x"a3c887ee",
   859 => x"49699749",
   860 => x"05a9c3c1",
   861 => x"a3c987dd",
   862 => x"49699749",
   863 => x"05a9c6c1",
   864 => x"a3ca87d1",
   865 => x"49699749",
   866 => x"05a9c7c1",
   867 => x"48c187c5",
   868 => x"c087e1c2",
   869 => x"87dcc248",
   870 => x"c087eafa",
   871 => x"f9f8c04c",
   872 => x"c049bf97",
   873 => x"87cf04a9",
   874 => x"c187fffa",
   875 => x"f9f8c084",
   876 => x"ac49bf97",
   877 => x"c087f106",
   878 => x"bf97f9f8",
   879 => x"f987cf02",
   880 => x"497087f8",
   881 => x"87c60299",
   882 => x"05a9ecc0",
   883 => x"4cc087f1",
   884 => x"7087e7f9",
   885 => x"87e2f94d",
   886 => x"f958a6c8",
   887 => x"4a7087dc",
   888 => x"a3c884c1",
   889 => x"49699749",
   890 => x"87c702ad",
   891 => x"05adffc0",
   892 => x"c987e7c0",
   893 => x"699749a3",
   894 => x"a966c449",
   895 => x"4887c702",
   896 => x"05a8ffc0",
   897 => x"a3ca87d4",
   898 => x"49699749",
   899 => x"87c602aa",
   900 => x"05aaffc0",
   901 => x"7ec187c4",
   902 => x"ecc087d0",
   903 => x"87c602ad",
   904 => x"05adfbc0",
   905 => x"4cc087c4",
   906 => x"026e7ec1",
   907 => x"f887e1fe",
   908 => x"487487ef",
   909 => x"ecfa8ef8",
   910 => x"5e0e0087",
   911 => x"0e5d5c5b",
   912 => x"c04b711e",
   913 => x"04ab4d4c",
   914 => x"c087e8c0",
   915 => x"751ed2f5",
   916 => x"87c4029d",
   917 => x"87c24ac0",
   918 => x"49724ac1",
   919 => x"c487e6ef",
   920 => x"c17e7086",
   921 => x"c2056e84",
   922 => x"c14c7387",
   923 => x"06ac7385",
   924 => x"6e87d8ff",
   925 => x"4d262648",
   926 => x"4b264c26",
   927 => x"5e0e4f26",
   928 => x"0e5d5c5b",
   929 => x"494c711e",
   930 => x"e7c291de",
   931 => x"85714dd9",
   932 => x"c1026d97",
   933 => x"e7c287dd",
   934 => x"744abfc4",
   935 => x"fe497282",
   936 => x"7e7087d8",
   937 => x"f3c0026e",
   938 => x"cce7c287",
   939 => x"cb4a6e4b",
   940 => x"f3c7ff49",
   941 => x"cb4b7487",
   942 => x"f2e0c193",
   943 => x"c083c483",
   944 => x"747bf7fb",
   945 => x"f4c6c149",
   946 => x"c27b7587",
   947 => x"bf97d8e7",
   948 => x"e7c21e49",
   949 => x"d9c149cc",
   950 => x"86c487f2",
   951 => x"c6c14974",
   952 => x"49c087db",
   953 => x"87fac7c1",
   954 => x"48c0e7c2",
   955 => x"49c178c0",
   956 => x"2687fddf",
   957 => x"4c87fffd",
   958 => x"6964616f",
   959 => x"2e2e676e",
   960 => x"5e0e002e",
   961 => x"710e5c5b",
   962 => x"e7c24a4b",
   963 => x"7282bfc4",
   964 => x"87e6fc49",
   965 => x"029c4c70",
   966 => x"eb4987c4",
   967 => x"e7c287ef",
   968 => x"78c048c4",
   969 => x"c7df49c1",
   970 => x"87ccfd87",
   971 => x"5c5b5e0e",
   972 => x"86f40e5d",
   973 => x"4dcedac2",
   974 => x"a6c44cc0",
   975 => x"c278c048",
   976 => x"49bfc4e7",
   977 => x"c106a9c0",
   978 => x"dac287c1",
   979 => x"029848ce",
   980 => x"c087f8c0",
   981 => x"c81ed2f5",
   982 => x"87c70266",
   983 => x"c048a6c4",
   984 => x"c487c578",
   985 => x"78c148a6",
   986 => x"eb4966c4",
   987 => x"86c487d7",
   988 => x"84c14d70",
   989 => x"c14866c4",
   990 => x"58a6c880",
   991 => x"bfc4e7c2",
   992 => x"c603ac49",
   993 => x"059d7587",
   994 => x"c087c8ff",
   995 => x"029d754c",
   996 => x"c087e0c3",
   997 => x"c81ed2f5",
   998 => x"87c70266",
   999 => x"c048a6cc",
  1000 => x"cc87c578",
  1001 => x"78c148a6",
  1002 => x"ea4966cc",
  1003 => x"86c487d7",
  1004 => x"026e7e70",
  1005 => x"6e87e9c2",
  1006 => x"9781cb49",
  1007 => x"99d04969",
  1008 => x"87d6c102",
  1009 => x"4ac2fcc0",
  1010 => x"91cb4974",
  1011 => x"81f2e0c1",
  1012 => x"81c87972",
  1013 => x"7451ffc3",
  1014 => x"c291de49",
  1015 => x"714dd9e7",
  1016 => x"97c1c285",
  1017 => x"49a5c17d",
  1018 => x"c251e0c0",
  1019 => x"bf97dee2",
  1020 => x"c187d202",
  1021 => x"4ba5c284",
  1022 => x"4adee2c2",
  1023 => x"c2ff49db",
  1024 => x"dbc187e6",
  1025 => x"49a5cd87",
  1026 => x"84c151c0",
  1027 => x"6e4ba5c2",
  1028 => x"ff49cb4a",
  1029 => x"c187d1c2",
  1030 => x"f9c087c6",
  1031 => x"49744afe",
  1032 => x"e0c191cb",
  1033 => x"797281f2",
  1034 => x"97dee2c2",
  1035 => x"87d802bf",
  1036 => x"91de4974",
  1037 => x"e7c284c1",
  1038 => x"83714bd9",
  1039 => x"4adee2c2",
  1040 => x"c1ff49dd",
  1041 => x"87d887e2",
  1042 => x"93de4b74",
  1043 => x"83d9e7c2",
  1044 => x"c049a3cb",
  1045 => x"7384c151",
  1046 => x"49cb4a6e",
  1047 => x"87c8c1ff",
  1048 => x"c14866c4",
  1049 => x"58a6c880",
  1050 => x"c003acc7",
  1051 => x"056e87c5",
  1052 => x"7487e0fc",
  1053 => x"f78ef448",
  1054 => x"731e87fc",
  1055 => x"494b711e",
  1056 => x"e0c191cb",
  1057 => x"a1c881f2",
  1058 => x"fad5c24a",
  1059 => x"c9501248",
  1060 => x"f8c04aa1",
  1061 => x"501248f9",
  1062 => x"e7c281ca",
  1063 => x"501148d8",
  1064 => x"97d8e7c2",
  1065 => x"c01e49bf",
  1066 => x"dfd2c149",
  1067 => x"c0e7c287",
  1068 => x"c178de48",
  1069 => x"87f8d849",
  1070 => x"87fef626",
  1071 => x"494a711e",
  1072 => x"e0c191cb",
  1073 => x"81c881f2",
  1074 => x"e7c24811",
  1075 => x"e7c258c4",
  1076 => x"78c048c4",
  1077 => x"d7d849c1",
  1078 => x"1e4f2687",
  1079 => x"c0c149c0",
  1080 => x"4f2687c0",
  1081 => x"0299711e",
  1082 => x"e2c187d2",
  1083 => x"50c048c7",
  1084 => x"c2c180f7",
  1085 => x"e0c140fc",
  1086 => x"87ce78e0",
  1087 => x"48c3e2c1",
  1088 => x"78c1e0c1",
  1089 => x"c3c180fc",
  1090 => x"4f2678db",
  1091 => x"5c5b5e0e",
  1092 => x"4a4c710e",
  1093 => x"e0c192cb",
  1094 => x"a2c882f2",
  1095 => x"4ba2c949",
  1096 => x"1e4b6b97",
  1097 => x"1e496997",
  1098 => x"491282ca",
  1099 => x"87fbeac0",
  1100 => x"fbd649c0",
  1101 => x"c0497487",
  1102 => x"f887c2fd",
  1103 => x"87f8f48e",
  1104 => x"711e731e",
  1105 => x"c3ff494b",
  1106 => x"fe497387",
  1107 => x"e9f487fe",
  1108 => x"1e731e87",
  1109 => x"a3c64b71",
  1110 => x"87dc024a",
  1111 => x"c0028ac1",
  1112 => x"028a87e4",
  1113 => x"8a87e8c1",
  1114 => x"87cac102",
  1115 => x"efc0028a",
  1116 => x"d9028a87",
  1117 => x"87e9c187",
  1118 => x"48c0e7c2",
  1119 => x"49c178df",
  1120 => x"c187edd5",
  1121 => x"49c787e6",
  1122 => x"c187f1fc",
  1123 => x"e7c287de",
  1124 => x"c102bfc4",
  1125 => x"c14887cb",
  1126 => x"c8e7c288",
  1127 => x"87c1c158",
  1128 => x"bfc8e7c2",
  1129 => x"87f9c002",
  1130 => x"bfc4e7c2",
  1131 => x"c280c148",
  1132 => x"c058c8e7",
  1133 => x"e7c287eb",
  1134 => x"c649bfc4",
  1135 => x"c8e7c289",
  1136 => x"a9b7c059",
  1137 => x"c287da03",
  1138 => x"c048c4e7",
  1139 => x"c287d278",
  1140 => x"02bfc8e7",
  1141 => x"e7c287cb",
  1142 => x"c648bfc4",
  1143 => x"c8e7c280",
  1144 => x"d449c058",
  1145 => x"497387ca",
  1146 => x"87d1fac0",
  1147 => x"0e87cbf2",
  1148 => x"0e5c5b5e",
  1149 => x"66cc4c71",
  1150 => x"cb4b741e",
  1151 => x"f2e0c193",
  1152 => x"4aa3c483",
  1153 => x"fafe496a",
  1154 => x"c1c187ee",
  1155 => x"a3c87bfa",
  1156 => x"5166d449",
  1157 => x"d849a3c9",
  1158 => x"a3ca5166",
  1159 => x"5166dc49",
  1160 => x"87d4f126",
  1161 => x"5c5b5e0e",
  1162 => x"d0ff0e5d",
  1163 => x"59a6d886",
  1164 => x"c048a6c8",
  1165 => x"c180fc78",
  1166 => x"c87866c4",
  1167 => x"c478c180",
  1168 => x"c278c180",
  1169 => x"c148c8e7",
  1170 => x"c0e7c278",
  1171 => x"486e7ebf",
  1172 => x"cb05a8de",
  1173 => x"87d4f387",
  1174 => x"a6cc4970",
  1175 => x"87f8d059",
  1176 => x"a8df486e",
  1177 => x"87eec105",
  1178 => x"4966c0c1",
  1179 => x"7e6981c4",
  1180 => x"48cddbc1",
  1181 => x"a1d0496e",
  1182 => x"7141204a",
  1183 => x"87f905aa",
  1184 => x"4afac1c1",
  1185 => x"0a66c0c1",
  1186 => x"c0c10a7a",
  1187 => x"81c94966",
  1188 => x"c0c151df",
  1189 => x"81ca4966",
  1190 => x"c151d3c1",
  1191 => x"cb4966c0",
  1192 => x"4ba1c481",
  1193 => x"6b48a6c4",
  1194 => x"721e7178",
  1195 => x"dddbc11e",
  1196 => x"4966cc48",
  1197 => x"204aa1d0",
  1198 => x"05aa7141",
  1199 => x"4a2687f9",
  1200 => x"79724926",
  1201 => x"df4aa1c9",
  1202 => x"c181ca52",
  1203 => x"a6c851d4",
  1204 => x"cf78c248",
  1205 => x"ece587c2",
  1206 => x"87cee687",
  1207 => x"7087dbe5",
  1208 => x"acfbc04c",
  1209 => x"87d0c102",
  1210 => x"c10566d4",
  1211 => x"1ec087c2",
  1212 => x"c11ec11e",
  1213 => x"c01ee5e2",
  1214 => x"87f3fb49",
  1215 => x"4a66d0c1",
  1216 => x"496a82c4",
  1217 => x"517481c7",
  1218 => x"1ed81ec1",
  1219 => x"81c8496a",
  1220 => x"d887ebe5",
  1221 => x"66c4c186",
  1222 => x"01a8c048",
  1223 => x"a6c887c7",
  1224 => x"ce78c148",
  1225 => x"66c4c187",
  1226 => x"c888c148",
  1227 => x"87c358a6",
  1228 => x"cc87f7e4",
  1229 => x"78c248a6",
  1230 => x"cd029c74",
  1231 => x"66c887d6",
  1232 => x"66c8c148",
  1233 => x"cbcd03a8",
  1234 => x"48a6d887",
  1235 => x"e9e378c0",
  1236 => x"c14c7087",
  1237 => x"c205acd0",
  1238 => x"66d887d6",
  1239 => x"87cde67e",
  1240 => x"a6dc4970",
  1241 => x"87d2e359",
  1242 => x"ecc04c70",
  1243 => x"eac105ac",
  1244 => x"4966c887",
  1245 => x"c0c191cb",
  1246 => x"a1c48166",
  1247 => x"c84d6a4a",
  1248 => x"66d84aa1",
  1249 => x"fcc2c152",
  1250 => x"87eee279",
  1251 => x"029c4c70",
  1252 => x"fbc087d8",
  1253 => x"87d202ac",
  1254 => x"dde25574",
  1255 => x"9c4c7087",
  1256 => x"c087c702",
  1257 => x"ff05acfb",
  1258 => x"e0c087ee",
  1259 => x"55c1c255",
  1260 => x"d47d97c0",
  1261 => x"a96e4966",
  1262 => x"c887db05",
  1263 => x"66c44866",
  1264 => x"87ca04a8",
  1265 => x"c14866c8",
  1266 => x"58a6cc80",
  1267 => x"66c487c8",
  1268 => x"c888c148",
  1269 => x"e1e158a6",
  1270 => x"c14c7087",
  1271 => x"c805acd0",
  1272 => x"4866d087",
  1273 => x"a6d480c1",
  1274 => x"acd0c158",
  1275 => x"87eafd02",
  1276 => x"d448a6dc",
  1277 => x"66d87866",
  1278 => x"a866dc48",
  1279 => x"87e6c905",
  1280 => x"48a6e0c0",
  1281 => x"c478f0c0",
  1282 => x"7866cc80",
  1283 => x"78c080c4",
  1284 => x"c048747e",
  1285 => x"f0c088fb",
  1286 => x"987058a6",
  1287 => x"87e1c802",
  1288 => x"c088cb48",
  1289 => x"7058a6f0",
  1290 => x"e9c00298",
  1291 => x"88c94887",
  1292 => x"58a6f0c0",
  1293 => x"c3029870",
  1294 => x"c44887e9",
  1295 => x"a6f0c088",
  1296 => x"02987058",
  1297 => x"c14887de",
  1298 => x"a6f0c088",
  1299 => x"02987058",
  1300 => x"c787d0c3",
  1301 => x"e0c087e5",
  1302 => x"78c048a6",
  1303 => x"c14866cc",
  1304 => x"58a6d080",
  1305 => x"87d2dfff",
  1306 => x"ecc04c70",
  1307 => x"87d702ac",
  1308 => x"0266e0c0",
  1309 => x"c087c7c0",
  1310 => x"c05ca6e4",
  1311 => x"487487c9",
  1312 => x"c088f0c0",
  1313 => x"c058a6e8",
  1314 => x"c002acec",
  1315 => x"deff87cd",
  1316 => x"4c7087e8",
  1317 => x"05acecc0",
  1318 => x"c087f3ff",
  1319 => x"d41e66e0",
  1320 => x"c01e4966",
  1321 => x"c11e66ec",
  1322 => x"d81ee5e2",
  1323 => x"fef44966",
  1324 => x"ca1ec087",
  1325 => x"66e0c01e",
  1326 => x"c191cb49",
  1327 => x"d88166d8",
  1328 => x"a1c448a6",
  1329 => x"bf66d878",
  1330 => x"f1deff49",
  1331 => x"c086d887",
  1332 => x"c106a8b7",
  1333 => x"1ec187c8",
  1334 => x"66c81ede",
  1335 => x"deff49bf",
  1336 => x"86c887dc",
  1337 => x"c0484970",
  1338 => x"e4c08808",
  1339 => x"b7c058a6",
  1340 => x"e9c006a8",
  1341 => x"66e0c087",
  1342 => x"a8b7dd48",
  1343 => x"6e87df03",
  1344 => x"e0c049bf",
  1345 => x"e0c08166",
  1346 => x"c1496651",
  1347 => x"81bf6e81",
  1348 => x"c051c1c2",
  1349 => x"c24966e0",
  1350 => x"81bf6e81",
  1351 => x"7ec151c0",
  1352 => x"ff87dec4",
  1353 => x"c087c6df",
  1354 => x"ff58a6e4",
  1355 => x"c087fede",
  1356 => x"c058a6e8",
  1357 => x"c005a8ec",
  1358 => x"e4c087cb",
  1359 => x"e0c048a6",
  1360 => x"c4c07866",
  1361 => x"f1dbff87",
  1362 => x"4966c887",
  1363 => x"c0c191cb",
  1364 => x"80714866",
  1365 => x"4a6e7e70",
  1366 => x"496e82c8",
  1367 => x"e0c081ca",
  1368 => x"e4c05166",
  1369 => x"81c14966",
  1370 => x"8966e0c0",
  1371 => x"307148c1",
  1372 => x"89c14970",
  1373 => x"c27a9771",
  1374 => x"49bff5ea",
  1375 => x"2966e0c0",
  1376 => x"484a6a97",
  1377 => x"f0c09871",
  1378 => x"496e58a6",
  1379 => x"4d6981c4",
  1380 => x"d84866dc",
  1381 => x"c002a866",
  1382 => x"a6d887c8",
  1383 => x"c078c048",
  1384 => x"a6d887c5",
  1385 => x"d878c148",
  1386 => x"e0c01e66",
  1387 => x"ff49751e",
  1388 => x"c887cbdb",
  1389 => x"c04c7086",
  1390 => x"c106acb7",
  1391 => x"857487d4",
  1392 => x"7449e0c0",
  1393 => x"c14b7589",
  1394 => x"714aeddb",
  1395 => x"87d8ebfe",
  1396 => x"e8c085c2",
  1397 => x"80c14866",
  1398 => x"58a6ecc0",
  1399 => x"4966ecc0",
  1400 => x"a97081c1",
  1401 => x"87c8c002",
  1402 => x"c048a6d8",
  1403 => x"87c5c078",
  1404 => x"c148a6d8",
  1405 => x"1e66d878",
  1406 => x"c049a4c2",
  1407 => x"887148e0",
  1408 => x"751e4970",
  1409 => x"f5d9ff49",
  1410 => x"c086c887",
  1411 => x"ff01a8b7",
  1412 => x"e8c087c0",
  1413 => x"d1c00266",
  1414 => x"c9496e87",
  1415 => x"66e8c081",
  1416 => x"c1486e51",
  1417 => x"c078ccc4",
  1418 => x"496e87cc",
  1419 => x"51c281c9",
  1420 => x"c5c1486e",
  1421 => x"7ec178c0",
  1422 => x"ff87c6c0",
  1423 => x"7087ebd8",
  1424 => x"c0026e4c",
  1425 => x"66c887f5",
  1426 => x"a866c448",
  1427 => x"87cbc004",
  1428 => x"c14866c8",
  1429 => x"58a6cc80",
  1430 => x"c487e0c0",
  1431 => x"88c14866",
  1432 => x"c058a6c8",
  1433 => x"c6c187d5",
  1434 => x"c8c005ac",
  1435 => x"4866cc87",
  1436 => x"a6d080c1",
  1437 => x"f1d7ff58",
  1438 => x"d04c7087",
  1439 => x"80c14866",
  1440 => x"7458a6d4",
  1441 => x"cbc0029c",
  1442 => x"4866c887",
  1443 => x"a866c8c1",
  1444 => x"87f5f204",
  1445 => x"87c9d7ff",
  1446 => x"c74866c8",
  1447 => x"e5c003a8",
  1448 => x"c8e7c287",
  1449 => x"c878c048",
  1450 => x"91cb4966",
  1451 => x"8166c0c1",
  1452 => x"6a4aa1c4",
  1453 => x"7952c04a",
  1454 => x"c14866c8",
  1455 => x"58a6cc80",
  1456 => x"ff04a8c7",
  1457 => x"d0ff87db",
  1458 => x"e9deff8e",
  1459 => x"616f4c87",
  1460 => x"65532064",
  1461 => x"6e697474",
  1462 => x"81207367",
  1463 => x"76615300",
  1464 => x"65532065",
  1465 => x"6e697474",
  1466 => x"81207367",
  1467 => x"00203a00",
  1468 => x"711e731e",
  1469 => x"c6029b4b",
  1470 => x"c4e7c287",
  1471 => x"c778c048",
  1472 => x"c4e7c21e",
  1473 => x"c11e49bf",
  1474 => x"c21ef2e0",
  1475 => x"49bfc0e7",
  1476 => x"cc87d1ec",
  1477 => x"c0e7c286",
  1478 => x"c7e749bf",
  1479 => x"029b7387",
  1480 => x"e0c187c8",
  1481 => x"e6c049f2",
  1482 => x"ddff87e5",
  1483 => x"731e87cc",
  1484 => x"c14bc01e",
  1485 => x"c049d9dd",
  1486 => x"c287fffa",
  1487 => x"c048fad5",
  1488 => x"d5e2c150",
  1489 => x"f4c049bf",
  1490 => x"987087d5",
  1491 => x"c187c405",
  1492 => x"734be5dd",
  1493 => x"e1dcff48",
  1494 => x"43495687",
  1495 => x"20203032",
  1496 => x"47464320",
  1497 => x"4d4f5200",
  1498 => x"616f6c20",
  1499 => x"676e6964",
  1500 => x"69616620",
  1501 => x"0064656c",
  1502 => x"87c8c81e",
  1503 => x"effd49c1",
  1504 => x"f6ecfe87",
  1505 => x"02987087",
  1506 => x"f5fe87cd",
  1507 => x"987087f3",
  1508 => x"c187c402",
  1509 => x"c087c24a",
  1510 => x"059a724a",
  1511 => x"1ec087ce",
  1512 => x"49ccdfc1",
  1513 => x"87f5f0c0",
  1514 => x"87fe86c4",
  1515 => x"87f4f7c0",
  1516 => x"dfc11ec0",
  1517 => x"f0c049d7",
  1518 => x"1ec087e3",
  1519 => x"7087effd",
  1520 => x"d8f0c049",
  1521 => x"87fbc387",
  1522 => x"4f268ef8",
  1523 => x"66204453",
  1524 => x"656c6961",
  1525 => x"42002e64",
  1526 => x"69746f6f",
  1527 => x"2e2e676e",
  1528 => x"c01e002e",
  1529 => x"fa87c4e8",
  1530 => x"1e4f2687",
  1531 => x"48c4e7c2",
  1532 => x"e7c278c0",
  1533 => x"78c048c0",
  1534 => x"e587fdfd",
  1535 => x"2648c087",
  1536 => x"2020204f",
  1537 => x"20202020",
  1538 => x"20202020",
  1539 => x"78452020",
  1540 => x"20207469",
  1541 => x"20202020",
  1542 => x"20202020",
  1543 => x"00812020",
  1544 => x"20202080",
  1545 => x"20202020",
  1546 => x"20202020",
  1547 => x"63614220",
  1548 => x"10bc006b",
  1549 => x"29d90000",
  1550 => x"00000000",
  1551 => x"0010bc00",
  1552 => x"0029f700",
  1553 => x"00000000",
  1554 => x"000010bc",
  1555 => x"00002a15",
  1556 => x"bc000000",
  1557 => x"33000010",
  1558 => x"0000002a",
  1559 => x"10bc0000",
  1560 => x"2a510000",
  1561 => x"00000000",
  1562 => x"0010bc00",
  1563 => x"002a6f00",
  1564 => x"00000000",
  1565 => x"000010bc",
  1566 => x"00002a8d",
  1567 => x"bc000000",
  1568 => x"00000010",
  1569 => x"00000000",
  1570 => x"11510000",
  1571 => x"00000000",
  1572 => x"00000000",
  1573 => x"00189900",
  1574 => x"43495600",
  1575 => x"20203032",
  1576 => x"4d4f5220",
  1577 => x"616f4c00",
  1578 => x"2e2a2064",
  1579 => x"f0fe1e00",
  1580 => x"cd78c048",
  1581 => x"26097909",
  1582 => x"fe1e1e4f",
  1583 => x"487ebff0",
  1584 => x"1e4f2626",
  1585 => x"c148f0fe",
  1586 => x"1e4f2678",
  1587 => x"c048f0fe",
  1588 => x"1e4f2678",
  1589 => x"52c04a71",
  1590 => x"0e4f2652",
  1591 => x"5d5c5b5e",
  1592 => x"7186f40e",
  1593 => x"7e6d974d",
  1594 => x"974ca5c1",
  1595 => x"a6c8486c",
  1596 => x"c4486e58",
  1597 => x"c505a866",
  1598 => x"c048ff87",
  1599 => x"caff87e6",
  1600 => x"49a5c287",
  1601 => x"714b6c97",
  1602 => x"6b974ba3",
  1603 => x"7e6c974b",
  1604 => x"80c1486e",
  1605 => x"c758a6c8",
  1606 => x"58a6cc98",
  1607 => x"fe7c9770",
  1608 => x"487387e1",
  1609 => x"4d268ef4",
  1610 => x"4b264c26",
  1611 => x"5e0e4f26",
  1612 => x"f40e5c5b",
  1613 => x"d84c7186",
  1614 => x"ffc34a66",
  1615 => x"4ba4c29a",
  1616 => x"73496c97",
  1617 => x"517249a1",
  1618 => x"6e7e6c97",
  1619 => x"c880c148",
  1620 => x"98c758a6",
  1621 => x"7058a6cc",
  1622 => x"ff8ef454",
  1623 => x"1e1e87ca",
  1624 => x"e087e8fd",
  1625 => x"c0494abf",
  1626 => x"0299c0e0",
  1627 => x"1e7287cb",
  1628 => x"49ebeac2",
  1629 => x"c487f7fe",
  1630 => x"87fdfc86",
  1631 => x"c2fd7e70",
  1632 => x"4f262687",
  1633 => x"ebeac21e",
  1634 => x"87c7fd49",
  1635 => x"49dee5c1",
  1636 => x"c587dafc",
  1637 => x"4f2687d9",
  1638 => x"5c5b5e0e",
  1639 => x"ebc20e5d",
  1640 => x"c14abfca",
  1641 => x"49bfece7",
  1642 => x"71bc724c",
  1643 => x"87dbfc4d",
  1644 => x"49744bc0",
  1645 => x"d50299d0",
  1646 => x"d0497587",
  1647 => x"c01e7199",
  1648 => x"feedc11e",
  1649 => x"1282734a",
  1650 => x"87e4c049",
  1651 => x"2cc186c8",
  1652 => x"abc8832d",
  1653 => x"87daff04",
  1654 => x"c187e8fb",
  1655 => x"c248ece7",
  1656 => x"78bfcaeb",
  1657 => x"4c264d26",
  1658 => x"4f264b26",
  1659 => x"00000000",
  1660 => x"48d0ff1e",
  1661 => x"ff78e1c8",
  1662 => x"78c548d4",
  1663 => x"c30266c4",
  1664 => x"78e0c387",
  1665 => x"c60266c8",
  1666 => x"48d4ff87",
  1667 => x"ff78f0c3",
  1668 => x"787148d4",
  1669 => x"c848d0ff",
  1670 => x"e0c078e1",
  1671 => x"0e4f2678",
  1672 => x"0e5c5b5e",
  1673 => x"eac24c71",
  1674 => x"eefa49eb",
  1675 => x"c04a7087",
  1676 => x"c204aab7",
  1677 => x"e0c387e3",
  1678 => x"87c905aa",
  1679 => x"48e2ebc1",
  1680 => x"d4c278c1",
  1681 => x"aaf0c387",
  1682 => x"c187c905",
  1683 => x"c148deeb",
  1684 => x"87f5c178",
  1685 => x"bfe2ebc1",
  1686 => x"7287c702",
  1687 => x"b3c0c24b",
  1688 => x"4b7287c2",
  1689 => x"d1059c74",
  1690 => x"deebc187",
  1691 => x"ebc11ebf",
  1692 => x"721ebfe2",
  1693 => x"87f8fd49",
  1694 => x"ebc186c8",
  1695 => x"c002bfde",
  1696 => x"497387e0",
  1697 => x"9129b7c4",
  1698 => x"81feecc1",
  1699 => x"9acf4a73",
  1700 => x"48c192c2",
  1701 => x"4a703072",
  1702 => x"4872baff",
  1703 => x"79709869",
  1704 => x"497387db",
  1705 => x"9129b7c4",
  1706 => x"81feecc1",
  1707 => x"9acf4a73",
  1708 => x"48c392c2",
  1709 => x"4a703072",
  1710 => x"70b06948",
  1711 => x"e2ebc179",
  1712 => x"c178c048",
  1713 => x"c048deeb",
  1714 => x"ebeac278",
  1715 => x"87cbf849",
  1716 => x"b7c04a70",
  1717 => x"ddfd03aa",
  1718 => x"fc48c087",
  1719 => x"000087c8",
  1720 => x"00000000",
  1721 => x"711e0000",
  1722 => x"f2fc494a",
  1723 => x"1e4f2687",
  1724 => x"49724ac0",
  1725 => x"ecc191c4",
  1726 => x"79c081fe",
  1727 => x"b7d082c1",
  1728 => x"87ee04aa",
  1729 => x"5e0e4f26",
  1730 => x"0e5d5c5b",
  1731 => x"faf64d71",
  1732 => x"c44a7587",
  1733 => x"c1922ab7",
  1734 => x"7582feec",
  1735 => x"c29ccf4c",
  1736 => x"4b496a94",
  1737 => x"9bc32b74",
  1738 => x"307448c2",
  1739 => x"bcff4c70",
  1740 => x"98714874",
  1741 => x"caf67a70",
  1742 => x"fa487387",
  1743 => x"000087e6",
  1744 => x"00000000",
  1745 => x"00000000",
  1746 => x"00000000",
  1747 => x"00000000",
  1748 => x"00000000",
  1749 => x"00000000",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"00000000",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"1e160000",
  1760 => x"362e2526",
  1761 => x"ff1e3e3d",
  1762 => x"e1c848d0",
  1763 => x"ff487178",
  1764 => x"c47808d4",
  1765 => x"d4ff4866",
  1766 => x"4f267808",
  1767 => x"c44a711e",
  1768 => x"e0c11e66",
  1769 => x"ddff49a2",
  1770 => x"4966c887",
  1771 => x"ff29b7c8",
  1772 => x"787148d4",
  1773 => x"c048d0ff",
  1774 => x"262678e0",
  1775 => x"d4ff1e4f",
  1776 => x"7affc34a",
  1777 => x"c848d0ff",
  1778 => x"7ade78e1",
  1779 => x"bff5eac2",
  1780 => x"c848497a",
  1781 => x"717a7028",
  1782 => x"7028d048",
  1783 => x"d848717a",
  1784 => x"ff7a7028",
  1785 => x"e0c048d0",
  1786 => x"0e4f2678",
  1787 => x"5d5c5b5e",
  1788 => x"c24c710e",
  1789 => x"4dbff5ea",
  1790 => x"d02b744b",
  1791 => x"83c19b66",
  1792 => x"04ab66d4",
  1793 => x"4bc087c2",
  1794 => x"66d04a74",
  1795 => x"ff317249",
  1796 => x"739975b9",
  1797 => x"70307248",
  1798 => x"b071484a",
  1799 => x"58f9eac2",
  1800 => x"2687dafe",
  1801 => x"264c264d",
  1802 => x"1e4f264b",
  1803 => x"c848d0ff",
  1804 => x"487178c9",
  1805 => x"7808d4ff",
  1806 => x"711e4f26",
  1807 => x"87eb494a",
  1808 => x"c848d0ff",
  1809 => x"1e4f2678",
  1810 => x"4b711e73",
  1811 => x"bfc5ebc2",
  1812 => x"c287c302",
  1813 => x"d0ff87eb",
  1814 => x"78c9c848",
  1815 => x"e0c04973",
  1816 => x"48d4ffb1",
  1817 => x"eac27871",
  1818 => x"78c048f9",
  1819 => x"c50266c8",
  1820 => x"49ffc387",
  1821 => x"49c087c2",
  1822 => x"59c1ebc2",
  1823 => x"c60266cc",
  1824 => x"d5d5c587",
  1825 => x"cf87c44a",
  1826 => x"c24affff",
  1827 => x"c25ac5eb",
  1828 => x"c148c5eb",
  1829 => x"2687c478",
  1830 => x"264c264d",
  1831 => x"0e4f264b",
  1832 => x"5d5c5b5e",
  1833 => x"c24a710e",
  1834 => x"4cbfc1eb",
  1835 => x"cb029a72",
  1836 => x"91c84987",
  1837 => x"4bfdf0c1",
  1838 => x"87c48371",
  1839 => x"4bfdf4c1",
  1840 => x"49134dc0",
  1841 => x"eac29974",
  1842 => x"ffb9bffd",
  1843 => x"787148d4",
  1844 => x"852cb7c1",
  1845 => x"04adb7c8",
  1846 => x"eac287e8",
  1847 => x"c848bff9",
  1848 => x"fdeac280",
  1849 => x"87effe58",
  1850 => x"711e731e",
  1851 => x"9a4a134b",
  1852 => x"7287cb02",
  1853 => x"87e7fe49",
  1854 => x"059a4a13",
  1855 => x"dafe87f5",
  1856 => x"eac21e87",
  1857 => x"c249bff9",
  1858 => x"c148f9ea",
  1859 => x"c0c478a1",
  1860 => x"db03a9b7",
  1861 => x"48d4ff87",
  1862 => x"bffdeac2",
  1863 => x"f9eac278",
  1864 => x"eac249bf",
  1865 => x"a1c148f9",
  1866 => x"b7c0c478",
  1867 => x"87e504a9",
  1868 => x"c848d0ff",
  1869 => x"c5ebc278",
  1870 => x"2678c048",
  1871 => x"0000004f",
  1872 => x"00000000",
  1873 => x"00000000",
  1874 => x"00005f5f",
  1875 => x"03030000",
  1876 => x"00030300",
  1877 => x"7f7f1400",
  1878 => x"147f7f14",
  1879 => x"2e240000",
  1880 => x"123a6b6b",
  1881 => x"366a4c00",
  1882 => x"32566c18",
  1883 => x"4f7e3000",
  1884 => x"683a7759",
  1885 => x"04000040",
  1886 => x"00000307",
  1887 => x"1c000000",
  1888 => x"0041633e",
  1889 => x"41000000",
  1890 => x"001c3e63",
  1891 => x"3e2a0800",
  1892 => x"2a3e1c1c",
  1893 => x"08080008",
  1894 => x"08083e3e",
  1895 => x"80000000",
  1896 => x"000060e0",
  1897 => x"08080000",
  1898 => x"08080808",
  1899 => x"00000000",
  1900 => x"00006060",
  1901 => x"30604000",
  1902 => x"03060c18",
  1903 => x"7f3e0001",
  1904 => x"3e7f4d59",
  1905 => x"06040000",
  1906 => x"00007f7f",
  1907 => x"63420000",
  1908 => x"464f5971",
  1909 => x"63220000",
  1910 => x"367f4949",
  1911 => x"161c1800",
  1912 => x"107f7f13",
  1913 => x"67270000",
  1914 => x"397d4545",
  1915 => x"7e3c0000",
  1916 => x"3079494b",
  1917 => x"01010000",
  1918 => x"070f7971",
  1919 => x"7f360000",
  1920 => x"367f4949",
  1921 => x"4f060000",
  1922 => x"1e3f6949",
  1923 => x"00000000",
  1924 => x"00006666",
  1925 => x"80000000",
  1926 => x"000066e6",
  1927 => x"08080000",
  1928 => x"22221414",
  1929 => x"14140000",
  1930 => x"14141414",
  1931 => x"22220000",
  1932 => x"08081414",
  1933 => x"03020000",
  1934 => x"060f5951",
  1935 => x"417f3e00",
  1936 => x"1e1f555d",
  1937 => x"7f7e0000",
  1938 => x"7e7f0909",
  1939 => x"7f7f0000",
  1940 => x"367f4949",
  1941 => x"3e1c0000",
  1942 => x"41414163",
  1943 => x"7f7f0000",
  1944 => x"1c3e6341",
  1945 => x"7f7f0000",
  1946 => x"41414949",
  1947 => x"7f7f0000",
  1948 => x"01010909",
  1949 => x"7f3e0000",
  1950 => x"7a7b4941",
  1951 => x"7f7f0000",
  1952 => x"7f7f0808",
  1953 => x"41000000",
  1954 => x"00417f7f",
  1955 => x"60200000",
  1956 => x"3f7f4040",
  1957 => x"087f7f00",
  1958 => x"4163361c",
  1959 => x"7f7f0000",
  1960 => x"40404040",
  1961 => x"067f7f00",
  1962 => x"7f7f060c",
  1963 => x"067f7f00",
  1964 => x"7f7f180c",
  1965 => x"7f3e0000",
  1966 => x"3e7f4141",
  1967 => x"7f7f0000",
  1968 => x"060f0909",
  1969 => x"417f3e00",
  1970 => x"407e7f61",
  1971 => x"7f7f0000",
  1972 => x"667f1909",
  1973 => x"6f260000",
  1974 => x"327b594d",
  1975 => x"01010000",
  1976 => x"01017f7f",
  1977 => x"7f3f0000",
  1978 => x"3f7f4040",
  1979 => x"3f0f0000",
  1980 => x"0f3f7070",
  1981 => x"307f7f00",
  1982 => x"7f7f3018",
  1983 => x"36634100",
  1984 => x"63361c1c",
  1985 => x"06030141",
  1986 => x"03067c7c",
  1987 => x"59716101",
  1988 => x"4143474d",
  1989 => x"7f000000",
  1990 => x"0041417f",
  1991 => x"06030100",
  1992 => x"6030180c",
  1993 => x"41000040",
  1994 => x"007f7f41",
  1995 => x"060c0800",
  1996 => x"080c0603",
  1997 => x"80808000",
  1998 => x"80808080",
  1999 => x"00000000",
  2000 => x"00040703",
  2001 => x"74200000",
  2002 => x"787c5454",
  2003 => x"7f7f0000",
  2004 => x"387c4444",
  2005 => x"7c380000",
  2006 => x"00444444",
  2007 => x"7c380000",
  2008 => x"7f7f4444",
  2009 => x"7c380000",
  2010 => x"185c5454",
  2011 => x"7e040000",
  2012 => x"0005057f",
  2013 => x"bc180000",
  2014 => x"7cfca4a4",
  2015 => x"7f7f0000",
  2016 => x"787c0404",
  2017 => x"00000000",
  2018 => x"00407d3d",
  2019 => x"80800000",
  2020 => x"007dfd80",
  2021 => x"7f7f0000",
  2022 => x"446c3810",
  2023 => x"00000000",
  2024 => x"00407f3f",
  2025 => x"0c7c7c00",
  2026 => x"787c0c18",
  2027 => x"7c7c0000",
  2028 => x"787c0404",
  2029 => x"7c380000",
  2030 => x"387c4444",
  2031 => x"fcfc0000",
  2032 => x"183c2424",
  2033 => x"3c180000",
  2034 => x"fcfc2424",
  2035 => x"7c7c0000",
  2036 => x"080c0404",
  2037 => x"5c480000",
  2038 => x"20745454",
  2039 => x"3f040000",
  2040 => x"0044447f",
  2041 => x"7c3c0000",
  2042 => x"7c7c4040",
  2043 => x"3c1c0000",
  2044 => x"1c3c6060",
  2045 => x"607c3c00",
  2046 => x"3c7c6030",
  2047 => x"386c4400",
  2048 => x"446c3810",
  2049 => x"bc1c0000",
  2050 => x"1c3c60e0",
  2051 => x"64440000",
  2052 => x"444c5c74",
  2053 => x"08080000",
  2054 => x"4141773e",
  2055 => x"00000000",
  2056 => x"00007f7f",
  2057 => x"41410000",
  2058 => x"08083e77",
  2059 => x"01010200",
  2060 => x"01020203",
  2061 => x"7f7f7f00",
  2062 => x"7f7f7f7f",
  2063 => x"1c080800",
  2064 => x"7f3e3e1c",
  2065 => x"3e7f7f7f",
  2066 => x"081c1c3e",
  2067 => x"18100008",
  2068 => x"10187c7c",
  2069 => x"30100000",
  2070 => x"10307c7c",
  2071 => x"60301000",
  2072 => x"061e7860",
  2073 => x"3c664200",
  2074 => x"42663c18",
  2075 => x"6a387800",
  2076 => x"386cc6c2",
  2077 => x"00006000",
  2078 => x"60000060",
  2079 => x"5b5e0e00",
  2080 => x"1e0e5d5c",
  2081 => x"ebc24c71",
  2082 => x"c04dbfd6",
  2083 => x"741ec04b",
  2084 => x"87c702ab",
  2085 => x"c048a6c4",
  2086 => x"c487c578",
  2087 => x"78c148a6",
  2088 => x"731e66c4",
  2089 => x"87dfee49",
  2090 => x"e0c086c8",
  2091 => x"87efef49",
  2092 => x"6a4aa5c4",
  2093 => x"87f0f049",
  2094 => x"cb87c6f1",
  2095 => x"c883c185",
  2096 => x"ff04abb7",
  2097 => x"262687c7",
  2098 => x"264c264d",
  2099 => x"1e4f264b",
  2100 => x"ebc24a71",
  2101 => x"ebc25ada",
  2102 => x"78c748da",
  2103 => x"87ddfe49",
  2104 => x"731e4f26",
  2105 => x"c04a711e",
  2106 => x"d303aab7",
  2107 => x"f2d0c287",
  2108 => x"87c405bf",
  2109 => x"87c24bc1",
  2110 => x"d0c24bc0",
  2111 => x"87c45bf6",
  2112 => x"5af6d0c2",
  2113 => x"bff2d0c2",
  2114 => x"c19ac14a",
  2115 => x"ec49a2c0",
  2116 => x"48fc87e8",
  2117 => x"bff2d0c2",
  2118 => x"87effe78",
  2119 => x"c44a711e",
  2120 => x"49721e66",
  2121 => x"2687f5e9",
  2122 => x"c21e4f26",
  2123 => x"49bff2d0",
  2124 => x"c287f3e6",
  2125 => x"e848ceeb",
  2126 => x"ebc278bf",
  2127 => x"bfec48ca",
  2128 => x"ceebc278",
  2129 => x"c3494abf",
  2130 => x"b7c899ff",
  2131 => x"7148722a",
  2132 => x"d6ebc2b0",
  2133 => x"0e4f2658",
  2134 => x"5d5c5b5e",
  2135 => x"ff4b710e",
  2136 => x"ebc287c8",
  2137 => x"50c048c9",
  2138 => x"d9e64973",
  2139 => x"4c497087",
  2140 => x"eecb9cc2",
  2141 => x"87c2cb49",
  2142 => x"c24d4970",
  2143 => x"bf97c9eb",
  2144 => x"87e2c105",
  2145 => x"c24966d0",
  2146 => x"99bfd2eb",
  2147 => x"d487d605",
  2148 => x"ebc24966",
  2149 => x"0599bfca",
  2150 => x"497387cb",
  2151 => x"7087e7e5",
  2152 => x"c1c10298",
  2153 => x"fe4cc187",
  2154 => x"497587c0",
  2155 => x"7087d7ca",
  2156 => x"87c60298",
  2157 => x"48c9ebc2",
  2158 => x"ebc250c1",
  2159 => x"05bf97c9",
  2160 => x"c287e3c0",
  2161 => x"49bfd2eb",
  2162 => x"059966d0",
  2163 => x"c287d6ff",
  2164 => x"49bfcaeb",
  2165 => x"059966d4",
  2166 => x"7387caff",
  2167 => x"87e6e449",
  2168 => x"fe059870",
  2169 => x"487487ff",
  2170 => x"0e87dcfb",
  2171 => x"5d5c5b5e",
  2172 => x"c086f40e",
  2173 => x"bfec4c4d",
  2174 => x"48a6c47e",
  2175 => x"bfd6ebc2",
  2176 => x"c01ec178",
  2177 => x"fd49c71e",
  2178 => x"86c887cd",
  2179 => x"cd029870",
  2180 => x"fb49ff87",
  2181 => x"dac187cc",
  2182 => x"87eae349",
  2183 => x"ebc24dc1",
  2184 => x"02bf97c9",
  2185 => x"d2cd87c3",
  2186 => x"ceebc287",
  2187 => x"d0c24bbf",
  2188 => x"c005bff2",
  2189 => x"fdc387e9",
  2190 => x"87cae349",
  2191 => x"e349fac3",
  2192 => x"497387c4",
  2193 => x"7199ffc3",
  2194 => x"fb49c01e",
  2195 => x"497387ce",
  2196 => x"7129b7c8",
  2197 => x"fb49c11e",
  2198 => x"86c887c2",
  2199 => x"c287f9c5",
  2200 => x"4bbfd2eb",
  2201 => x"87dd029b",
  2202 => x"bfeed0c2",
  2203 => x"87d6c749",
  2204 => x"c4059870",
  2205 => x"d24bc087",
  2206 => x"49e0c287",
  2207 => x"c287fbc6",
  2208 => x"c658f2d0",
  2209 => x"eed0c287",
  2210 => x"7378c048",
  2211 => x"0599c249",
  2212 => x"ebc387cd",
  2213 => x"87eee149",
  2214 => x"99c24970",
  2215 => x"fb87c202",
  2216 => x"c149734c",
  2217 => x"87cd0599",
  2218 => x"e149f4c3",
  2219 => x"497087d8",
  2220 => x"c20299c2",
  2221 => x"734cfa87",
  2222 => x"0599c849",
  2223 => x"f5c387cd",
  2224 => x"87c2e149",
  2225 => x"99c24970",
  2226 => x"c287d402",
  2227 => x"02bfdaeb",
  2228 => x"c14887c9",
  2229 => x"deebc288",
  2230 => x"ff87c258",
  2231 => x"734dc14c",
  2232 => x"0599c449",
  2233 => x"f2c387cd",
  2234 => x"87dae049",
  2235 => x"99c24970",
  2236 => x"c287db02",
  2237 => x"7ebfdaeb",
  2238 => x"a8b7c748",
  2239 => x"6e87cb03",
  2240 => x"c280c148",
  2241 => x"c058deeb",
  2242 => x"4cfe87c2",
  2243 => x"fdc34dc1",
  2244 => x"f1dfff49",
  2245 => x"c2497087",
  2246 => x"87d50299",
  2247 => x"bfdaebc2",
  2248 => x"87c9c002",
  2249 => x"48daebc2",
  2250 => x"c2c078c0",
  2251 => x"c14cfd87",
  2252 => x"49fac34d",
  2253 => x"87cedfff",
  2254 => x"99c24970",
  2255 => x"c287d902",
  2256 => x"48bfdaeb",
  2257 => x"03a8b7c7",
  2258 => x"c287c9c0",
  2259 => x"c748daeb",
  2260 => x"87c2c078",
  2261 => x"4dc14cfc",
  2262 => x"03acb7c0",
  2263 => x"c487d1c0",
  2264 => x"d8c14a66",
  2265 => x"c0026a82",
  2266 => x"4b6a87c6",
  2267 => x"0f734974",
  2268 => x"f0c31ec0",
  2269 => x"49dac11e",
  2270 => x"c887dcf7",
  2271 => x"02987086",
  2272 => x"c887e2c0",
  2273 => x"ebc248a6",
  2274 => x"c878bfda",
  2275 => x"91cb4966",
  2276 => x"714866c4",
  2277 => x"6e7e7080",
  2278 => x"c8c002bf",
  2279 => x"4bbf6e87",
  2280 => x"734966c8",
  2281 => x"029d750f",
  2282 => x"c287c8c0",
  2283 => x"49bfdaeb",
  2284 => x"c287caf3",
  2285 => x"02bff6d0",
  2286 => x"4987ddc0",
  2287 => x"7087c7c2",
  2288 => x"d3c00298",
  2289 => x"daebc287",
  2290 => x"f0f249bf",
  2291 => x"f449c087",
  2292 => x"d0c287d0",
  2293 => x"78c048f6",
  2294 => x"eaf38ef4",
  2295 => x"5b5e0e87",
  2296 => x"1e0e5d5c",
  2297 => x"ebc24c71",
  2298 => x"c149bfd6",
  2299 => x"c14da1cd",
  2300 => x"7e6981d1",
  2301 => x"cf029c74",
  2302 => x"4ba5c487",
  2303 => x"ebc27b74",
  2304 => x"f349bfd6",
  2305 => x"7b6e87c9",
  2306 => x"c4059c74",
  2307 => x"c24bc087",
  2308 => x"734bc187",
  2309 => x"87caf349",
  2310 => x"c70266d4",
  2311 => x"87da4987",
  2312 => x"87c24a70",
  2313 => x"d0c24ac0",
  2314 => x"f2265afa",
  2315 => x"000087d9",
  2316 => x"00000000",
  2317 => x"00000000",
  2318 => x"711e0000",
  2319 => x"bfc8ff4a",
  2320 => x"48a17249",
  2321 => x"ff1e4f26",
  2322 => x"fe89bfc8",
  2323 => x"c0c0c0c0",
  2324 => x"c401a9c0",
  2325 => x"c24ac087",
  2326 => x"724ac187",
  2327 => x"0e4f2648",
  2328 => x"5d5c5b5e",
  2329 => x"7e711e0e",
  2330 => x"6e4bd4ff",
  2331 => x"deebc21e",
  2332 => x"d8cffe49",
  2333 => x"7086c487",
  2334 => x"c3029d4d",
  2335 => x"ebc287c3",
  2336 => x"6e4cbfe6",
  2337 => x"d0e2fe49",
  2338 => x"48d0ff87",
  2339 => x"c178c5c8",
  2340 => x"4ac07bd6",
  2341 => x"82c17b15",
  2342 => x"aab7e0c0",
  2343 => x"ff87f504",
  2344 => x"78c448d0",
  2345 => x"c178c5c8",
  2346 => x"7bc17bd3",
  2347 => x"9c7478c4",
  2348 => x"87fcc102",
  2349 => x"7ecedac2",
  2350 => x"8c4dc0c8",
  2351 => x"03acb7c0",
  2352 => x"c0c887c6",
  2353 => x"4cc04da4",
  2354 => x"97ffe6c2",
  2355 => x"99d049bf",
  2356 => x"c087d202",
  2357 => x"deebc21e",
  2358 => x"ccd1fe49",
  2359 => x"7086c487",
  2360 => x"efc04a49",
  2361 => x"cedac287",
  2362 => x"deebc21e",
  2363 => x"f8d0fe49",
  2364 => x"7086c487",
  2365 => x"d0ff4a49",
  2366 => x"78c5c848",
  2367 => x"6e7bd4c1",
  2368 => x"6e7bbf97",
  2369 => x"7080c148",
  2370 => x"058dc17e",
  2371 => x"ff87f0ff",
  2372 => x"78c448d0",
  2373 => x"c5059a72",
  2374 => x"c048c087",
  2375 => x"1ec187e5",
  2376 => x"49deebc2",
  2377 => x"87e0cefe",
  2378 => x"9c7486c4",
  2379 => x"87c4fe05",
  2380 => x"c848d0ff",
  2381 => x"d3c178c5",
  2382 => x"c47bc07b",
  2383 => x"c248c178",
  2384 => x"2648c087",
  2385 => x"4c264d26",
  2386 => x"4f264b26",
  2387 => x"711e731e",
  2388 => x"0266c84a",
  2389 => x"c14b87ce",
  2390 => x"ce028bd3",
  2391 => x"028bc187",
  2392 => x"87d387d0",
  2393 => x"f6fb4972",
  2394 => x"7287cc87",
  2395 => x"87cac249",
  2396 => x"497287c5",
  2397 => x"ff87f6c2",
  2398 => x"1e0087ce",
  2399 => x"bfe2d9c2",
  2400 => x"c2b9c149",
  2401 => x"ff59e6d9",
  2402 => x"ffc348d4",
  2403 => x"48d0ff78",
  2404 => x"ff78e1c8",
  2405 => x"78c148d4",
  2406 => x"787131c4",
  2407 => x"c048d0ff",
  2408 => x"4f2678e0",
  2409 => x"fdd6c21e",
  2410 => x"deebc21e",
  2411 => x"dccafe49",
  2412 => x"7086c487",
  2413 => x"87c30298",
  2414 => x"2687c0ff",
  2415 => x"4b35314f",
  2416 => x"20205a48",
  2417 => x"47464320",
  2418 => x"4a711e00",
  2419 => x"c249a2c4",
  2420 => x"6a48f5ea",
  2421 => x"c1496978",
  2422 => x"e6d9c2b9",
  2423 => x"87dbfe59",
  2424 => x"87d9d7ff",
  2425 => x"4f2648c1",
  2426 => x"c44a711e",
  2427 => x"eac249a2",
  2428 => x"c27abff5",
  2429 => x"79bfe2d9",
  2430 => x"711e4f26",
  2431 => x"ebc21e4a",
  2432 => x"c9fe49de",
  2433 => x"86c487c7",
  2434 => x"dc029870",
  2435 => x"cedac287",
  2436 => x"deebc21e",
  2437 => x"d0ccfe49",
  2438 => x"7086c487",
  2439 => x"87c90298",
  2440 => x"49cedac2",
  2441 => x"c287e2fe",
  2442 => x"2648c087",
  2443 => x"4a711e4f",
  2444 => x"deebc21e",
  2445 => x"d4c8fe49",
  2446 => x"7086c487",
  2447 => x"87de0298",
  2448 => x"49cedac2",
  2449 => x"c287e1fe",
  2450 => x"c21eceda",
  2451 => x"fe49deeb",
  2452 => x"c487d9cc",
  2453 => x"02987086",
  2454 => x"48c187c4",
  2455 => x"48c087c2",
  2456 => x"00004f26",
  2457 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
