library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"446c3810",
     1 => x"bc1c0000",
     2 => x"1c3c60e0",
     3 => x"64440000",
     4 => x"444c5c74",
     5 => x"08080000",
     6 => x"4141773e",
     7 => x"00000000",
     8 => x"00007f7f",
     9 => x"41410000",
    10 => x"08083e77",
    11 => x"01010200",
    12 => x"01020203",
    13 => x"7f7f7f00",
    14 => x"7f7f7f7f",
    15 => x"1c080800",
    16 => x"7f3e3e1c",
    17 => x"3e7f7f7f",
    18 => x"081c1c3e",
    19 => x"18100008",
    20 => x"10187c7c",
    21 => x"30100000",
    22 => x"10307c7c",
    23 => x"60301000",
    24 => x"061e7860",
    25 => x"3c664200",
    26 => x"42663c18",
    27 => x"6a387800",
    28 => x"386cc6c2",
    29 => x"00006000",
    30 => x"60000060",
    31 => x"5b5e0e00",
    32 => x"1e0e5d5c",
    33 => x"ebc24c71",
    34 => x"c04dbfd6",
    35 => x"741ec04b",
    36 => x"87c702ab",
    37 => x"c048a6c4",
    38 => x"c487c578",
    39 => x"78c148a6",
    40 => x"731e66c4",
    41 => x"87dfee49",
    42 => x"e0c086c8",
    43 => x"87efef49",
    44 => x"6a4aa5c4",
    45 => x"87f0f049",
    46 => x"cb87c6f1",
    47 => x"c883c185",
    48 => x"ff04abb7",
    49 => x"262687c7",
    50 => x"264c264d",
    51 => x"1e4f264b",
    52 => x"ebc24a71",
    53 => x"ebc25ada",
    54 => x"78c748da",
    55 => x"87ddfe49",
    56 => x"731e4f26",
    57 => x"c04a711e",
    58 => x"d303aab7",
    59 => x"f2d0c287",
    60 => x"87c405bf",
    61 => x"87c24bc1",
    62 => x"d0c24bc0",
    63 => x"87c45bf6",
    64 => x"5af6d0c2",
    65 => x"bff2d0c2",
    66 => x"c19ac14a",
    67 => x"ec49a2c0",
    68 => x"48fc87e8",
    69 => x"bff2d0c2",
    70 => x"87effe78",
    71 => x"c44a711e",
    72 => x"49721e66",
    73 => x"2687f5e9",
    74 => x"c21e4f26",
    75 => x"49bff2d0",
    76 => x"c287f3e6",
    77 => x"e848ceeb",
    78 => x"ebc278bf",
    79 => x"bfec48ca",
    80 => x"ceebc278",
    81 => x"c3494abf",
    82 => x"b7c899ff",
    83 => x"7148722a",
    84 => x"d6ebc2b0",
    85 => x"0e4f2658",
    86 => x"5d5c5b5e",
    87 => x"ff4b710e",
    88 => x"ebc287c8",
    89 => x"50c048c9",
    90 => x"d9e64973",
    91 => x"4c497087",
    92 => x"eecb9cc2",
    93 => x"87c2cb49",
    94 => x"c24d4970",
    95 => x"bf97c9eb",
    96 => x"87e2c105",
    97 => x"c24966d0",
    98 => x"99bfd2eb",
    99 => x"d487d605",
   100 => x"ebc24966",
   101 => x"0599bfca",
   102 => x"497387cb",
   103 => x"7087e7e5",
   104 => x"c1c10298",
   105 => x"fe4cc187",
   106 => x"497587c0",
   107 => x"7087d7ca",
   108 => x"87c60298",
   109 => x"48c9ebc2",
   110 => x"ebc250c1",
   111 => x"05bf97c9",
   112 => x"c287e3c0",
   113 => x"49bfd2eb",
   114 => x"059966d0",
   115 => x"c287d6ff",
   116 => x"49bfcaeb",
   117 => x"059966d4",
   118 => x"7387caff",
   119 => x"87e6e449",
   120 => x"fe059870",
   121 => x"487487ff",
   122 => x"0e87dcfb",
   123 => x"5d5c5b5e",
   124 => x"c086f40e",
   125 => x"bfec4c4d",
   126 => x"48a6c47e",
   127 => x"bfd6ebc2",
   128 => x"c01ec178",
   129 => x"fd49c71e",
   130 => x"86c887cd",
   131 => x"cd029870",
   132 => x"fb49ff87",
   133 => x"dac187cc",
   134 => x"87eae349",
   135 => x"ebc24dc1",
   136 => x"02bf97c9",
   137 => x"d2cd87c3",
   138 => x"ceebc287",
   139 => x"d0c24bbf",
   140 => x"c005bff2",
   141 => x"fdc387e9",
   142 => x"87cae349",
   143 => x"e349fac3",
   144 => x"497387c4",
   145 => x"7199ffc3",
   146 => x"fb49c01e",
   147 => x"497387ce",
   148 => x"7129b7c8",
   149 => x"fb49c11e",
   150 => x"86c887c2",
   151 => x"c287f9c5",
   152 => x"4bbfd2eb",
   153 => x"87dd029b",
   154 => x"bfeed0c2",
   155 => x"87d6c749",
   156 => x"c4059870",
   157 => x"d24bc087",
   158 => x"49e0c287",
   159 => x"c287fbc6",
   160 => x"c658f2d0",
   161 => x"eed0c287",
   162 => x"7378c048",
   163 => x"0599c249",
   164 => x"ebc387cd",
   165 => x"87eee149",
   166 => x"99c24970",
   167 => x"fb87c202",
   168 => x"c149734c",
   169 => x"87cd0599",
   170 => x"e149f4c3",
   171 => x"497087d8",
   172 => x"c20299c2",
   173 => x"734cfa87",
   174 => x"0599c849",
   175 => x"f5c387cd",
   176 => x"87c2e149",
   177 => x"99c24970",
   178 => x"c287d402",
   179 => x"02bfdaeb",
   180 => x"c14887c9",
   181 => x"deebc288",
   182 => x"ff87c258",
   183 => x"734dc14c",
   184 => x"0599c449",
   185 => x"f2c387cd",
   186 => x"87dae049",
   187 => x"99c24970",
   188 => x"c287db02",
   189 => x"7ebfdaeb",
   190 => x"a8b7c748",
   191 => x"6e87cb03",
   192 => x"c280c148",
   193 => x"c058deeb",
   194 => x"4cfe87c2",
   195 => x"fdc34dc1",
   196 => x"f1dfff49",
   197 => x"c2497087",
   198 => x"87d50299",
   199 => x"bfdaebc2",
   200 => x"87c9c002",
   201 => x"48daebc2",
   202 => x"c2c078c0",
   203 => x"c14cfd87",
   204 => x"49fac34d",
   205 => x"87cedfff",
   206 => x"99c24970",
   207 => x"c287d902",
   208 => x"48bfdaeb",
   209 => x"03a8b7c7",
   210 => x"c287c9c0",
   211 => x"c748daeb",
   212 => x"87c2c078",
   213 => x"4dc14cfc",
   214 => x"03acb7c0",
   215 => x"c487d1c0",
   216 => x"d8c14a66",
   217 => x"c0026a82",
   218 => x"4b6a87c6",
   219 => x"0f734974",
   220 => x"f0c31ec0",
   221 => x"49dac11e",
   222 => x"c887dcf7",
   223 => x"02987086",
   224 => x"c887e2c0",
   225 => x"ebc248a6",
   226 => x"c878bfda",
   227 => x"91cb4966",
   228 => x"714866c4",
   229 => x"6e7e7080",
   230 => x"c8c002bf",
   231 => x"4bbf6e87",
   232 => x"734966c8",
   233 => x"029d750f",
   234 => x"c287c8c0",
   235 => x"49bfdaeb",
   236 => x"c287caf3",
   237 => x"02bff6d0",
   238 => x"4987ddc0",
   239 => x"7087c7c2",
   240 => x"d3c00298",
   241 => x"daebc287",
   242 => x"f0f249bf",
   243 => x"f449c087",
   244 => x"d0c287d0",
   245 => x"78c048f6",
   246 => x"eaf38ef4",
   247 => x"5b5e0e87",
   248 => x"1e0e5d5c",
   249 => x"ebc24c71",
   250 => x"c149bfd6",
   251 => x"c14da1cd",
   252 => x"7e6981d1",
   253 => x"cf029c74",
   254 => x"4ba5c487",
   255 => x"ebc27b74",
   256 => x"f349bfd6",
   257 => x"7b6e87c9",
   258 => x"c4059c74",
   259 => x"c24bc087",
   260 => x"734bc187",
   261 => x"87caf349",
   262 => x"c70266d4",
   263 => x"87da4987",
   264 => x"87c24a70",
   265 => x"d0c24ac0",
   266 => x"f2265afa",
   267 => x"000087d9",
   268 => x"00000000",
   269 => x"00000000",
   270 => x"711e0000",
   271 => x"bfc8ff4a",
   272 => x"48a17249",
   273 => x"ff1e4f26",
   274 => x"fe89bfc8",
   275 => x"c0c0c0c0",
   276 => x"c401a9c0",
   277 => x"c24ac087",
   278 => x"724ac187",
   279 => x"0e4f2648",
   280 => x"5d5c5b5e",
   281 => x"7e711e0e",
   282 => x"6e4bd4ff",
   283 => x"deebc21e",
   284 => x"d8cffe49",
   285 => x"7086c487",
   286 => x"c3029d4d",
   287 => x"ebc287c3",
   288 => x"6e4cbfe6",
   289 => x"d0e2fe49",
   290 => x"48d0ff87",
   291 => x"c178c5c8",
   292 => x"4ac07bd6",
   293 => x"82c17b15",
   294 => x"aab7e0c0",
   295 => x"ff87f504",
   296 => x"78c448d0",
   297 => x"c178c5c8",
   298 => x"7bc17bd3",
   299 => x"9c7478c4",
   300 => x"87fcc102",
   301 => x"7ecedac2",
   302 => x"8c4dc0c8",
   303 => x"03acb7c0",
   304 => x"c0c887c6",
   305 => x"4cc04da4",
   306 => x"97ffe6c2",
   307 => x"99d049bf",
   308 => x"c087d202",
   309 => x"deebc21e",
   310 => x"ccd1fe49",
   311 => x"7086c487",
   312 => x"efc04a49",
   313 => x"cedac287",
   314 => x"deebc21e",
   315 => x"f8d0fe49",
   316 => x"7086c487",
   317 => x"d0ff4a49",
   318 => x"78c5c848",
   319 => x"6e7bd4c1",
   320 => x"6e7bbf97",
   321 => x"7080c148",
   322 => x"058dc17e",
   323 => x"ff87f0ff",
   324 => x"78c448d0",
   325 => x"c5059a72",
   326 => x"c048c087",
   327 => x"1ec187e5",
   328 => x"49deebc2",
   329 => x"87e0cefe",
   330 => x"9c7486c4",
   331 => x"87c4fe05",
   332 => x"c848d0ff",
   333 => x"d3c178c5",
   334 => x"c47bc07b",
   335 => x"c248c178",
   336 => x"2648c087",
   337 => x"4c264d26",
   338 => x"4f264b26",
   339 => x"711e731e",
   340 => x"0266c84a",
   341 => x"c14b87ce",
   342 => x"ce028bd3",
   343 => x"028bc187",
   344 => x"87d387d0",
   345 => x"f6fb4972",
   346 => x"7287cc87",
   347 => x"87cac249",
   348 => x"497287c5",
   349 => x"ff87f6c2",
   350 => x"1e0087ce",
   351 => x"bfe2d9c2",
   352 => x"c2b9c149",
   353 => x"ff59e6d9",
   354 => x"ffc348d4",
   355 => x"48d0ff78",
   356 => x"ff78e1c8",
   357 => x"78c148d4",
   358 => x"787131c4",
   359 => x"c048d0ff",
   360 => x"4f2678e0",
   361 => x"fdd6c21e",
   362 => x"deebc21e",
   363 => x"dccafe49",
   364 => x"7086c487",
   365 => x"87c30298",
   366 => x"2687c0ff",
   367 => x"4b35314f",
   368 => x"20205a48",
   369 => x"47464320",
   370 => x"4a711e00",
   371 => x"c249a2c4",
   372 => x"6a48f5ea",
   373 => x"c1496978",
   374 => x"e6d9c2b9",
   375 => x"87dbfe59",
   376 => x"87d9d7ff",
   377 => x"4f2648c1",
   378 => x"c44a711e",
   379 => x"eac249a2",
   380 => x"c27abff5",
   381 => x"79bfe2d9",
   382 => x"711e4f26",
   383 => x"ebc21e4a",
   384 => x"c9fe49de",
   385 => x"86c487c7",
   386 => x"dc029870",
   387 => x"cedac287",
   388 => x"deebc21e",
   389 => x"d0ccfe49",
   390 => x"7086c487",
   391 => x"87c90298",
   392 => x"49cedac2",
   393 => x"c287e2fe",
   394 => x"2648c087",
   395 => x"4a711e4f",
   396 => x"deebc21e",
   397 => x"d4c8fe49",
   398 => x"7086c487",
   399 => x"87de0298",
   400 => x"49cedac2",
   401 => x"c287e1fe",
   402 => x"c21eceda",
   403 => x"fe49deeb",
   404 => x"c487d9cc",
   405 => x"02987086",
   406 => x"48c187c4",
   407 => x"48c087c2",
   408 => x"00004f26",
   409 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
